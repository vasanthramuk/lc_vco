magic
tech sky130A
timestamp 1670733274
<< pwell >>
rect -148 -1673 148 1673
<< nmos >>
rect -50 1028 50 1568
rect -50 379 50 919
rect -50 -270 50 270
rect -50 -919 50 -379
rect -50 -1568 50 -1028
<< ndiff >>
rect -79 1562 -50 1568
rect -79 1034 -73 1562
rect -56 1034 -50 1562
rect -79 1028 -50 1034
rect 50 1562 79 1568
rect 50 1034 56 1562
rect 73 1034 79 1562
rect 50 1028 79 1034
rect -79 913 -50 919
rect -79 385 -73 913
rect -56 385 -50 913
rect -79 379 -50 385
rect 50 913 79 919
rect 50 385 56 913
rect 73 385 79 913
rect 50 379 79 385
rect -79 264 -50 270
rect -79 -264 -73 264
rect -56 -264 -50 264
rect -79 -270 -50 -264
rect 50 264 79 270
rect 50 -264 56 264
rect 73 -264 79 264
rect 50 -270 79 -264
rect -79 -385 -50 -379
rect -79 -913 -73 -385
rect -56 -913 -50 -385
rect -79 -919 -50 -913
rect 50 -385 79 -379
rect 50 -913 56 -385
rect 73 -913 79 -385
rect 50 -919 79 -913
rect -79 -1034 -50 -1028
rect -79 -1562 -73 -1034
rect -56 -1562 -50 -1034
rect -79 -1568 -50 -1562
rect 50 -1034 79 -1028
rect 50 -1562 56 -1034
rect 73 -1562 79 -1034
rect 50 -1568 79 -1562
<< ndiffc >>
rect -73 1034 -56 1562
rect 56 1034 73 1562
rect -73 385 -56 913
rect 56 385 73 913
rect -73 -264 -56 264
rect 56 -264 73 264
rect -73 -913 -56 -385
rect 56 -913 73 -385
rect -73 -1562 -56 -1034
rect 56 -1562 73 -1034
<< psubdiff >>
rect -130 1638 -82 1655
rect 82 1638 130 1655
rect -130 1607 -113 1638
rect 113 1607 130 1638
rect -130 -1638 -113 -1607
rect 113 -1638 130 -1607
rect -130 -1655 -82 -1638
rect 82 -1655 130 -1638
<< psubdiffcont >>
rect -82 1638 82 1655
rect -130 -1607 -113 1607
rect 113 -1607 130 1607
rect -82 -1655 82 -1638
<< poly >>
rect -50 1604 50 1612
rect -50 1587 -42 1604
rect 42 1587 50 1604
rect -50 1568 50 1587
rect -50 1009 50 1028
rect -50 992 -42 1009
rect 42 992 50 1009
rect -50 984 50 992
rect -50 955 50 963
rect -50 938 -42 955
rect 42 938 50 955
rect -50 919 50 938
rect -50 360 50 379
rect -50 343 -42 360
rect 42 343 50 360
rect -50 335 50 343
rect -50 306 50 314
rect -50 289 -42 306
rect 42 289 50 306
rect -50 270 50 289
rect -50 -289 50 -270
rect -50 -306 -42 -289
rect 42 -306 50 -289
rect -50 -314 50 -306
rect -50 -343 50 -335
rect -50 -360 -42 -343
rect 42 -360 50 -343
rect -50 -379 50 -360
rect -50 -938 50 -919
rect -50 -955 -42 -938
rect 42 -955 50 -938
rect -50 -963 50 -955
rect -50 -992 50 -984
rect -50 -1009 -42 -992
rect 42 -1009 50 -992
rect -50 -1028 50 -1009
rect -50 -1587 50 -1568
rect -50 -1604 -42 -1587
rect 42 -1604 50 -1587
rect -50 -1612 50 -1604
<< polycont >>
rect -42 1587 42 1604
rect -42 992 42 1009
rect -42 938 42 955
rect -42 343 42 360
rect -42 289 42 306
rect -42 -306 42 -289
rect -42 -360 42 -343
rect -42 -955 42 -938
rect -42 -1009 42 -992
rect -42 -1604 42 -1587
<< locali >>
rect -130 1638 -82 1655
rect 82 1638 130 1655
rect -130 1607 -113 1638
rect 113 1607 130 1638
rect -50 1587 -42 1604
rect 42 1587 50 1604
rect -73 1562 -56 1570
rect -73 1026 -56 1034
rect 56 1562 73 1570
rect 56 1026 73 1034
rect -50 992 -42 1009
rect 42 992 50 1009
rect -50 938 -42 955
rect 42 938 50 955
rect -73 913 -56 921
rect -73 377 -56 385
rect 56 913 73 921
rect 56 377 73 385
rect -50 343 -42 360
rect 42 343 50 360
rect -50 289 -42 306
rect 42 289 50 306
rect -73 264 -56 272
rect -73 -272 -56 -264
rect 56 264 73 272
rect 56 -272 73 -264
rect -50 -306 -42 -289
rect 42 -306 50 -289
rect -50 -360 -42 -343
rect 42 -360 50 -343
rect -73 -385 -56 -377
rect -73 -921 -56 -913
rect 56 -385 73 -377
rect 56 -921 73 -913
rect -50 -955 -42 -938
rect 42 -955 50 -938
rect -50 -1009 -42 -992
rect 42 -1009 50 -992
rect -73 -1034 -56 -1026
rect -73 -1570 -56 -1562
rect 56 -1034 73 -1026
rect 56 -1570 73 -1562
rect -50 -1604 -42 -1587
rect 42 -1604 50 -1587
rect -130 -1638 -113 -1607
rect 113 -1638 130 -1607
rect -130 -1655 -82 -1638
rect 82 -1655 130 -1638
<< viali >>
rect -42 1587 42 1604
rect -73 1034 -56 1562
rect 56 1034 73 1562
rect -42 992 42 1009
rect -42 938 42 955
rect -73 385 -56 913
rect 56 385 73 913
rect -42 343 42 360
rect -42 289 42 306
rect -73 -264 -56 264
rect 56 -264 73 264
rect -42 -306 42 -289
rect -42 -360 42 -343
rect -73 -913 -56 -385
rect 56 -913 73 -385
rect -42 -955 42 -938
rect -42 -1009 42 -992
rect -73 -1562 -56 -1034
rect 56 -1562 73 -1034
rect -42 -1604 42 -1587
<< metal1 >>
rect -48 1604 48 1607
rect -48 1587 -42 1604
rect 42 1587 48 1604
rect -48 1584 48 1587
rect -76 1562 -53 1568
rect -76 1034 -73 1562
rect -56 1034 -53 1562
rect -76 1028 -53 1034
rect 53 1562 76 1568
rect 53 1034 56 1562
rect 73 1034 76 1562
rect 53 1028 76 1034
rect -48 1009 48 1012
rect -48 992 -42 1009
rect 42 992 48 1009
rect -48 989 48 992
rect -48 955 48 958
rect -48 938 -42 955
rect 42 938 48 955
rect -48 935 48 938
rect -76 913 -53 919
rect -76 385 -73 913
rect -56 385 -53 913
rect -76 379 -53 385
rect 53 913 76 919
rect 53 385 56 913
rect 73 385 76 913
rect 53 379 76 385
rect -48 360 48 363
rect -48 343 -42 360
rect 42 343 48 360
rect -48 340 48 343
rect -48 306 48 309
rect -48 289 -42 306
rect 42 289 48 306
rect -48 286 48 289
rect -76 264 -53 270
rect -76 -264 -73 264
rect -56 -264 -53 264
rect -76 -270 -53 -264
rect 53 264 76 270
rect 53 -264 56 264
rect 73 -264 76 264
rect 53 -270 76 -264
rect -48 -289 48 -286
rect -48 -306 -42 -289
rect 42 -306 48 -289
rect -48 -309 48 -306
rect -48 -343 48 -340
rect -48 -360 -42 -343
rect 42 -360 48 -343
rect -48 -363 48 -360
rect -76 -385 -53 -379
rect -76 -913 -73 -385
rect -56 -913 -53 -385
rect -76 -919 -53 -913
rect 53 -385 76 -379
rect 53 -913 56 -385
rect 73 -913 76 -385
rect 53 -919 76 -913
rect -48 -938 48 -935
rect -48 -955 -42 -938
rect 42 -955 48 -938
rect -48 -958 48 -955
rect -48 -992 48 -989
rect -48 -1009 -42 -992
rect 42 -1009 48 -992
rect -48 -1012 48 -1009
rect -76 -1034 -53 -1028
rect -76 -1562 -73 -1034
rect -56 -1562 -53 -1034
rect -76 -1568 -53 -1562
rect 53 -1034 76 -1028
rect 53 -1562 56 -1034
rect 73 -1562 76 -1034
rect 53 -1568 76 -1562
rect -48 -1587 48 -1584
rect -48 -1604 -42 -1587
rect 42 -1604 48 -1587
rect -48 -1607 48 -1604
<< properties >>
string FIXED_BBOX -121 -1646 121 1646
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.4 l 1 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
