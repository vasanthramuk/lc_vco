* SPICE3 file created from sonamutha.ext - technology: sky130A

X0 vp curgate curgate vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X1 vp curgate curgate vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X2 vp m3_5645_4434# m2_2622_5196# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3 vp m2_2622_5196# m3_5645_4434# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4 m3_5645_4434# m2_2622_5196# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5 vp m2_2622_5196# m3_5645_4434# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 m2_2622_5196# m3_5645_4434# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7 vp m3_5645_4434# m2_2622_5196# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8 m3_5645_4434# m2_2622_5196# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 m2_2622_5196# m3_5645_4434# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10 m2_2622_5196# m1_2705_3336# vp sky130_fd_pr__cap_var_lvt w=1e+07u l=500000u
X11 m3_5645_4434# m1_2705_3336# vp sky130_fd_pr__cap_var_lvt w=1e+07u l=500000u
X12 VDD m2_2622_5196# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X13 VDD m3_5645_4434# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X14 VDD m2_2622_5196# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X15 VDD m3_5645_4434# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X16 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X17 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X18 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X19 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X20 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
C0 m3_5645_4434# m1_2705_3336# 2.46fF
C1 VDD m2_2622_5196# 88.19fF
C2 m3_5645_4434# m2_2622_5196# 5.31fF
C3 VDD m3_5645_4434# 88.21fF
C4 m1_2705_3336# m2_2622_5196# 2.40fF
C5 curgate vp 6.22fF **FLOATING
C6 VDD vp 8.20fF **FLOATING
C7 m1_2705_3336# vp 9.14fF **FLOATING
C8 m3_5645_4434# vp 28.28fF **FLOATING
C9 m2_2622_5196# vp 29.78fF **FLOATING
C10 sky130_fd_pr__nfet_01v8_TPE47J_0/w_n1018_n1448# vp 7.16fF **FLOATING
