magic
tech sky130A
magscale 1 2
timestamp 1671534598
<< nwell >>
rect 1532 4640 4222 4906
rect 1532 2104 1962 4640
rect 3888 2104 4222 4640
rect 1532 1826 4222 2104
<< pwell >>
rect -55 6699 537 9497
rect -53 -53 539 6639
rect 1962 2104 3888 4640
<< nmos >>
rect 141 8207 341 9287
rect 141 6909 341 7989
rect 143 5349 343 6429
rect 143 4051 343 5131
rect 143 2753 343 3833
rect 143 1455 343 2535
rect 143 157 343 1237
rect 2397 3481 2597 4281
rect 2655 3481 2855 4281
rect 2913 3481 3113 4281
rect 3171 3481 3371 4281
rect 2397 2463 2597 3263
rect 2655 2463 2855 3263
rect 2913 2463 3113 3263
rect 3171 2463 3371 3263
<< ndiff >>
rect 83 9275 141 9287
rect 83 8219 95 9275
rect 129 8219 141 9275
rect 83 8207 141 8219
rect 341 9275 399 9287
rect 341 8219 353 9275
rect 387 8219 399 9275
rect 341 8207 399 8219
rect 83 7977 141 7989
rect 83 6921 95 7977
rect 129 6921 141 7977
rect 83 6909 141 6921
rect 341 7977 399 7989
rect 341 6921 353 7977
rect 387 6921 399 7977
rect 341 6909 399 6921
rect 85 6417 143 6429
rect 85 5361 97 6417
rect 131 5361 143 6417
rect 85 5349 143 5361
rect 343 6417 401 6429
rect 343 5361 355 6417
rect 389 5361 401 6417
rect 343 5349 401 5361
rect 85 5119 143 5131
rect 85 4063 97 5119
rect 131 4063 143 5119
rect 85 4051 143 4063
rect 343 5119 401 5131
rect 343 4063 355 5119
rect 389 4063 401 5119
rect 343 4051 401 4063
rect 85 3821 143 3833
rect 85 2765 97 3821
rect 131 2765 143 3821
rect 85 2753 143 2765
rect 343 3821 401 3833
rect 343 2765 355 3821
rect 389 2765 401 3821
rect 343 2753 401 2765
rect 85 2523 143 2535
rect 85 1467 97 2523
rect 131 1467 143 2523
rect 85 1455 143 1467
rect 343 2523 401 2535
rect 343 1467 355 2523
rect 389 1467 401 2523
rect 343 1455 401 1467
rect 85 1225 143 1237
rect 85 169 97 1225
rect 131 169 143 1225
rect 85 157 143 169
rect 343 1225 401 1237
rect 343 169 355 1225
rect 389 169 401 1225
rect 343 157 401 169
rect 2339 4269 2397 4281
rect 2339 3493 2351 4269
rect 2385 3493 2397 4269
rect 2339 3481 2397 3493
rect 2597 4269 2655 4281
rect 2597 3493 2609 4269
rect 2643 3493 2655 4269
rect 2597 3481 2655 3493
rect 2855 4269 2913 4281
rect 2855 3493 2867 4269
rect 2901 3493 2913 4269
rect 2855 3481 2913 3493
rect 3113 4269 3171 4281
rect 3113 3493 3125 4269
rect 3159 3493 3171 4269
rect 3113 3481 3171 3493
rect 3371 4269 3429 4281
rect 3371 3493 3383 4269
rect 3417 3493 3429 4269
rect 3371 3481 3429 3493
rect 2339 3251 2397 3263
rect 2339 2475 2351 3251
rect 2385 2475 2397 3251
rect 2339 2463 2397 2475
rect 2597 3251 2655 3263
rect 2597 2475 2609 3251
rect 2643 2475 2655 3251
rect 2597 2463 2655 2475
rect 2855 3251 2913 3263
rect 2855 2475 2867 3251
rect 2901 2475 2913 3251
rect 2855 2463 2913 2475
rect 3113 3251 3171 3263
rect 3113 2475 3125 3251
rect 3159 2475 3171 3251
rect 3113 2463 3171 2475
rect 3371 3251 3429 3263
rect 3371 2475 3383 3251
rect 3417 2475 3429 3251
rect 3371 2463 3429 2475
<< ndiffc >>
rect 95 8219 129 9275
rect 353 8219 387 9275
rect 95 6921 129 7977
rect 353 6921 387 7977
rect 97 5361 131 6417
rect 355 5361 389 6417
rect 97 4063 131 5119
rect 355 4063 389 5119
rect 97 2765 131 3821
rect 355 2765 389 3821
rect 97 1467 131 2523
rect 355 1467 389 2523
rect 97 169 131 1225
rect 355 169 389 1225
rect 2351 3493 2385 4269
rect 2609 3493 2643 4269
rect 2867 3493 2901 4269
rect 3125 3493 3159 4269
rect 3383 3493 3417 4269
rect 2351 2475 2385 3251
rect 2609 2475 2643 3251
rect 2867 2475 2901 3251
rect 3125 2475 3159 3251
rect 3383 2475 3417 3251
<< psubdiff >>
rect -19 9427 77 9461
rect 405 9427 501 9461
rect -19 9365 15 9427
rect -919 8014 -802 8039
rect -919 7967 -887 8014
rect -829 7967 -802 8014
rect -919 7943 -802 7967
rect 467 9365 501 9427
rect -19 6769 15 6831
rect 467 6769 501 6831
rect -19 6735 77 6769
rect 405 6735 501 6769
rect -17 6569 79 6603
rect 407 6569 503 6603
rect -17 6507 17 6569
rect 469 6507 503 6569
rect -17 17 17 79
rect 2237 4421 2333 4455
rect 3435 4421 3531 4455
rect 2237 4359 2271 4421
rect 3497 4359 3531 4421
rect 2237 2323 2271 2385
rect 3497 2323 3531 2385
rect 2237 2289 2333 2323
rect 3435 2289 3531 2323
rect 469 17 503 79
rect -17 -17 79 17
rect 407 -17 503 17
<< nsubdiff >>
rect 3980 4822 4148 4848
rect 1646 4806 4148 4822
rect 1646 4690 1670 4806
rect 4086 4706 4148 4806
rect 1648 1926 1670 4690
rect 1794 4690 4002 4706
rect 1794 2044 1816 4690
rect 3978 2044 4002 4690
rect 1794 2024 4002 2044
rect 4084 4694 4148 4706
rect 4084 2024 4108 4694
rect 4086 1926 4108 2024
rect 1648 1902 4108 1926
<< psubdiffcont >>
rect 77 9427 405 9461
rect -887 7967 -829 8014
rect -19 6831 15 9365
rect 467 6831 501 9365
rect 77 6735 405 6769
rect 79 6569 407 6603
rect -17 79 17 6507
rect 469 79 503 6507
rect 2333 4421 3435 4455
rect 2237 2385 2271 4359
rect 3497 2385 3531 4359
rect 2333 2289 3435 2323
rect 79 -17 407 17
<< nsubdiffcont >>
rect 1670 4706 4086 4806
rect 1670 2024 1794 4706
rect 4002 2024 4084 4706
rect 1670 1926 4086 2024
<< poly >>
rect 141 9359 341 9375
rect 141 9325 157 9359
rect 325 9325 341 9359
rect 141 9287 341 9325
rect 141 8136 341 8207
rect 141 8061 258 8136
rect 316 8061 341 8136
rect 141 7989 341 8061
rect 141 6871 341 6909
rect 141 6837 157 6871
rect 325 6837 341 6871
rect 141 6821 341 6837
rect 143 6501 343 6517
rect 143 6467 159 6501
rect 327 6467 343 6501
rect 143 6429 343 6467
rect 143 5131 343 5349
rect 143 3833 343 4051
rect 143 2535 343 2753
rect 143 1237 343 1455
rect 143 69 343 157
rect 2397 4353 2597 4369
rect 2397 4319 2413 4353
rect 2581 4319 2597 4353
rect 2397 4281 2597 4319
rect 2655 4353 2855 4369
rect 2655 4319 2671 4353
rect 2839 4319 2855 4353
rect 2655 4281 2855 4319
rect 2913 4353 3113 4369
rect 2913 4319 2929 4353
rect 3097 4319 3113 4353
rect 2913 4281 3113 4319
rect 3171 4353 3371 4369
rect 3171 4319 3187 4353
rect 3355 4319 3371 4353
rect 3171 4281 3371 4319
rect 2397 3443 2597 3481
rect 2397 3409 2413 3443
rect 2581 3409 2597 3443
rect 2397 3393 2597 3409
rect 2655 3443 2855 3481
rect 2655 3409 2671 3443
rect 2839 3409 2855 3443
rect 2655 3393 2855 3409
rect 2913 3443 3113 3481
rect 2913 3409 2929 3443
rect 3097 3409 3113 3443
rect 2913 3393 3113 3409
rect 3171 3443 3371 3481
rect 3171 3409 3187 3443
rect 3355 3409 3371 3443
rect 3171 3393 3371 3409
rect 2397 3335 2597 3351
rect 2397 3301 2413 3335
rect 2581 3301 2597 3335
rect 2397 3263 2597 3301
rect 2655 3335 2855 3351
rect 2655 3301 2671 3335
rect 2839 3301 2855 3335
rect 2655 3263 2855 3301
rect 2913 3335 3113 3351
rect 2913 3301 2929 3335
rect 3097 3301 3113 3335
rect 2913 3263 3113 3301
rect 3171 3335 3371 3351
rect 3171 3301 3187 3335
rect 3355 3301 3371 3335
rect 3171 3263 3371 3301
rect 2397 2425 2597 2463
rect 2397 2391 2413 2425
rect 2581 2391 2597 2425
rect 2397 2375 2597 2391
rect 2655 2425 2855 2463
rect 2655 2391 2671 2425
rect 2839 2391 2855 2425
rect 2655 2375 2855 2391
rect 2913 2425 3113 2463
rect 2913 2391 2929 2425
rect 3097 2391 3113 2425
rect 2913 2375 3113 2391
rect 3171 2425 3371 2463
rect 3171 2391 3187 2425
rect 3355 2391 3371 2425
rect 3171 2375 3371 2391
<< polycont >>
rect 157 9325 325 9359
rect 258 8061 316 8136
rect 157 6837 325 6871
rect 159 6467 327 6501
rect 2413 4319 2581 4353
rect 2671 4319 2839 4353
rect 2929 4319 3097 4353
rect 3187 4319 3355 4353
rect 2413 3409 2581 3443
rect 2671 3409 2839 3443
rect 2929 3409 3097 3443
rect 3187 3409 3355 3443
rect 2413 3301 2581 3335
rect 2671 3301 2839 3335
rect 2929 3301 3097 3335
rect 3187 3301 3355 3335
rect 2413 2391 2581 2425
rect 2671 2391 2839 2425
rect 2929 2391 3097 2425
rect 3187 2391 3355 2425
<< locali >>
rect -19 9427 77 9461
rect 405 9427 501 9461
rect -19 9365 15 9427
rect -910 8014 -807 8037
rect -910 7967 -887 8014
rect -829 7967 -807 8014
rect -218 7988 -19 8214
rect -910 7948 -807 7967
rect 467 9365 501 9427
rect 141 9325 157 9359
rect 325 9325 341 9359
rect 95 9275 129 9291
rect 95 8214 129 8219
rect 15 7984 129 8214
rect 353 9275 387 9291
rect 353 8156 387 8219
rect 244 8136 387 8156
rect 244 8061 258 8136
rect 316 8061 387 8136
rect 244 8039 387 8061
rect 95 7977 129 7984
rect 95 6905 129 6921
rect 353 7977 387 8039
rect 353 6905 387 6921
rect 141 6837 157 6871
rect 325 6837 341 6871
rect -19 6769 15 6831
rect 467 6769 501 6831
rect -19 6735 77 6769
rect 405 6735 501 6769
rect -17 6569 79 6603
rect 407 6569 503 6603
rect -17 6507 17 6569
rect -370 2768 -17 3820
rect 469 6507 503 6569
rect 143 6467 159 6501
rect 327 6467 343 6501
rect 97 6417 131 6433
rect 97 5119 131 5361
rect 97 3821 131 4063
rect 17 2766 97 3820
rect 355 6417 389 6433
rect 355 5119 389 5361
rect 355 3821 389 4063
rect 354 3056 355 3494
rect 97 2523 131 2765
rect 97 1225 131 1467
rect 97 153 131 169
rect 355 2523 389 2765
rect 355 1225 389 1467
rect 355 153 389 169
rect -17 17 17 79
rect 1630 4806 4122 4836
rect 1630 2190 1670 4806
rect 4086 4706 4122 4806
rect 1311 1926 1670 2190
rect 1794 4702 4002 4706
rect 1794 2066 1880 4702
rect 2237 4421 2333 4455
rect 3435 4421 3531 4455
rect 2237 4359 2271 4421
rect 2230 4234 2237 4240
rect 3497 4359 3531 4421
rect 2397 4319 2413 4353
rect 2581 4319 2597 4353
rect 2655 4319 2671 4353
rect 2839 4319 2855 4353
rect 2913 4319 2929 4353
rect 3097 4319 3113 4353
rect 3171 4319 3187 4353
rect 3355 4319 3371 4353
rect 2351 4269 2385 4285
rect 2271 4234 2282 4240
rect 2609 4269 2643 4285
rect 2230 4118 2236 4234
rect 2272 4118 2282 4234
rect 2230 4112 2237 4118
rect 2228 2620 2237 2626
rect 2271 4112 2282 4118
rect 2351 3477 2385 3493
rect 2867 4269 2901 4285
rect 3125 4269 3159 4285
rect 2609 3477 2643 3493
rect 3383 4269 3417 4285
rect 3490 4236 3497 4240
rect 3531 4236 3540 4240
rect 3490 4118 3496 4236
rect 3532 4118 3540 4236
rect 2867 3477 2901 3493
rect 3125 3477 3159 3493
rect 3490 4112 3497 4118
rect 3383 3477 3417 3493
rect 2397 3409 2413 3443
rect 2581 3409 2597 3443
rect 2655 3409 2671 3443
rect 2839 3409 2855 3443
rect 2913 3409 2929 3443
rect 3097 3409 3113 3443
rect 3171 3409 3187 3443
rect 3355 3409 3371 3443
rect 2397 3301 2413 3335
rect 2581 3301 2597 3335
rect 2655 3301 2671 3335
rect 2839 3301 2855 3335
rect 2913 3301 2929 3335
rect 3097 3301 3113 3335
rect 3171 3301 3187 3335
rect 3355 3301 3371 3335
rect 2351 3251 2385 3267
rect 2271 2620 2282 2626
rect 2609 3251 2643 3267
rect 2867 3251 2901 3267
rect 2228 2504 2236 2620
rect 2272 2504 2282 2620
rect 2228 2496 2237 2504
rect 2271 2496 2282 2504
rect 2351 2459 2385 2475
rect 3125 3251 3159 3267
rect 3383 3251 3417 3267
rect 2609 2459 2643 2475
rect 2867 2459 2901 2475
rect 3487 2619 3497 2622
rect 3531 4112 3540 4118
rect 3531 2619 3539 2622
rect 3125 2459 3159 2475
rect 3487 2503 3496 2619
rect 3532 2503 3539 2619
rect 3487 2495 3497 2503
rect 3383 2459 3417 2475
rect 2397 2391 2413 2425
rect 2581 2391 2597 2425
rect 2655 2391 2671 2425
rect 2839 2391 2855 2425
rect 2913 2391 2929 2425
rect 3097 2391 3113 2425
rect 3171 2391 3187 2425
rect 3355 2391 3371 2425
rect 2237 2323 2271 2385
rect 3531 2495 3539 2503
rect 3497 2323 3531 2385
rect 2237 2289 2333 2323
rect 3435 2289 3531 2323
rect 3964 2066 4002 4702
rect 1794 2024 4002 2066
rect 4084 2066 4122 4706
rect 4084 2024 4124 2066
rect 4086 1926 4124 2024
rect 1311 1901 4124 1926
rect 1630 1878 4124 1901
rect 1630 1874 1880 1878
rect 469 17 503 79
rect -17 -17 79 17
rect 407 -17 503 17
<< viali >>
rect 157 9325 325 9359
rect 157 6837 325 6871
rect 159 6467 327 6501
rect 355 2765 389 3821
rect 2413 4319 2581 4353
rect 2671 4319 2839 4353
rect 2929 4319 3097 4353
rect 3187 4319 3355 4353
rect 2236 4118 2237 4234
rect 2237 4118 2271 4234
rect 2271 4118 2272 4234
rect 2350 4118 2351 4234
rect 2351 4118 2385 4234
rect 2385 4118 2386 4234
rect 2866 4116 2867 4234
rect 2867 4116 2901 4234
rect 2901 4116 2902 4234
rect 2610 3638 2643 3752
rect 2643 3638 2644 3752
rect 3382 4116 3383 4234
rect 3383 4116 3417 4234
rect 3417 4116 3418 4234
rect 3496 4118 3497 4236
rect 3497 4118 3531 4236
rect 3531 4118 3532 4236
rect 3124 3638 3125 3752
rect 3125 3638 3158 3752
rect 2413 3409 2581 3443
rect 2671 3409 2839 3443
rect 2929 3409 3097 3443
rect 3187 3409 3355 3443
rect 2413 3301 2581 3335
rect 2671 3301 2839 3335
rect 2929 3301 3097 3335
rect 3187 3301 3355 3335
rect 2606 2994 2609 3110
rect 2609 2994 2643 3110
rect 2643 2994 2646 3110
rect 2236 2504 2237 2620
rect 2237 2504 2271 2620
rect 2271 2504 2272 2620
rect 2350 2504 2351 2620
rect 2351 2504 2385 2620
rect 2385 2504 2386 2620
rect 3122 2998 3125 3112
rect 3125 2998 3159 3112
rect 3159 2998 3162 3112
rect 2866 2504 2867 2620
rect 2867 2504 2901 2620
rect 2901 2504 2902 2620
rect 3382 2504 3383 2620
rect 3383 2504 3417 2620
rect 3417 2504 3418 2620
rect 3496 2503 3497 2619
rect 3497 2503 3531 2619
rect 3531 2503 3532 2619
rect 2413 2391 2581 2425
rect 2671 2391 2839 2425
rect 2929 2391 3097 2425
rect 3187 2391 3355 2425
<< metal1 >>
rect 145 9359 337 9365
rect 145 9325 157 9359
rect 325 9325 337 9359
rect 145 9319 337 9325
rect 145 6871 337 6877
rect 145 6837 157 6871
rect 325 6837 337 6871
rect 145 6831 337 6837
rect 146 6507 337 6831
rect 146 6501 339 6507
rect 146 6467 159 6501
rect 327 6467 339 6501
rect 146 6462 339 6467
rect 147 6461 339 6462
rect 2401 4353 2593 4359
rect 2401 4319 2413 4353
rect 2581 4319 2593 4353
rect 2401 4313 2593 4319
rect 2659 4353 2851 4359
rect 2659 4319 2671 4353
rect 2839 4319 2851 4353
rect 2659 4313 2851 4319
rect 2917 4353 3109 4359
rect 2917 4319 2929 4353
rect 3097 4319 3109 4353
rect 2917 4313 3109 4319
rect 3175 4353 3367 4359
rect 3175 4319 3187 4353
rect 3355 4319 3367 4353
rect 3175 4313 3367 4319
rect 1200 4246 2427 4248
rect 1200 4236 3548 4246
rect 1200 4234 3496 4236
rect 1200 4118 2236 4234
rect 2272 4118 2350 4234
rect 2386 4118 2866 4234
rect 1200 4116 2866 4118
rect 2902 4116 3382 4234
rect 3418 4118 3496 4234
rect 3532 4118 3548 4236
rect 3418 4116 3548 4118
rect 1200 4100 3548 4116
rect 1200 4099 2427 4100
rect 582 3836 930 3840
rect 1200 3836 1474 4099
rect 340 3821 1014 3836
rect 340 2765 355 3821
rect 389 3384 1014 3821
rect 1124 3384 1479 3836
rect 2594 3752 3178 3762
rect 2594 3638 2610 3752
rect 2644 3690 3124 3752
rect 2644 3638 2684 3690
rect 2594 3634 2684 3638
rect 2836 3638 3124 3690
rect 3158 3638 3178 3752
rect 2836 3634 3178 3638
rect 2594 3624 3178 3634
rect 2918 3449 3110 3450
rect 2401 3448 2593 3449
rect 2659 3448 2851 3449
rect 2917 3448 3110 3449
rect 3175 3448 3367 3449
rect 2401 3446 3367 3448
rect 2401 3443 2924 3446
rect 3106 3443 3367 3446
rect 2401 3409 2413 3443
rect 2581 3409 2671 3443
rect 2839 3409 2924 3443
rect 3106 3409 3187 3443
rect 3355 3409 3367 3443
rect 2401 3404 2924 3409
rect 2401 3403 2593 3404
rect 2659 3403 2851 3404
rect 2917 3403 2924 3404
rect 2918 3392 2924 3403
rect 3106 3404 3367 3409
rect 3106 3392 3110 3404
rect 3175 3403 3367 3404
rect 2918 3386 3110 3392
rect 389 3212 1479 3384
rect 2658 3356 2856 3360
rect 2401 3340 2593 3341
rect 2658 3340 2664 3356
rect 2401 3335 2664 3340
rect 2850 3340 2856 3356
rect 2917 3340 3109 3341
rect 3175 3340 3367 3341
rect 2850 3335 3367 3340
rect 2401 3301 2413 3335
rect 2581 3301 2664 3335
rect 2850 3301 2929 3335
rect 3097 3301 3187 3335
rect 3355 3301 3367 3335
rect 2401 3298 2664 3301
rect 2850 3298 3367 3301
rect 2401 3295 2593 3298
rect 2658 3296 2856 3298
rect 2659 3295 2851 3296
rect 2917 3295 3109 3298
rect 3175 3295 3367 3298
rect 389 2765 1014 3212
rect 340 2750 1014 2765
rect 872 2749 1014 2750
rect 1124 2749 1479 3212
rect 2590 3122 3184 3128
rect 2590 3110 2946 3122
rect 2590 2994 2606 3110
rect 2646 3066 2946 3110
rect 3098 3112 3184 3122
rect 3098 3066 3122 3112
rect 2646 2998 3122 3066
rect 3162 2998 3184 3112
rect 2646 2994 3184 2998
rect 2590 2982 3184 2994
rect 1198 2630 1479 2749
rect 2340 2631 3446 2632
rect 2340 2630 3530 2631
rect 1198 2620 3548 2630
rect 1198 2504 2236 2620
rect 2272 2504 2350 2620
rect 2386 2504 2866 2620
rect 2902 2504 3382 2620
rect 3418 2619 3548 2620
rect 3418 2504 3496 2619
rect 1198 2503 3496 2504
rect 3532 2503 3548 2619
rect 1198 2482 3548 2503
rect 3399 2481 3548 2482
rect 3480 2480 3548 2481
rect 2401 2430 2593 2431
rect 2659 2430 2851 2431
rect 2917 2430 3109 2431
rect 3175 2430 3367 2431
rect 2401 2425 3367 2430
rect 2401 2391 2413 2425
rect 2581 2391 2671 2425
rect 2839 2391 2929 2425
rect 3097 2391 3187 2425
rect 3355 2391 3367 2425
rect 2401 2386 3367 2391
rect 2401 2385 2593 2386
rect 2659 2385 2851 2386
rect 2917 2385 3109 2386
rect 3175 2385 3367 2386
<< via1 >>
rect 2684 3634 2836 3690
rect 2924 3443 3106 3446
rect 2924 3409 2929 3443
rect 2929 3409 3097 3443
rect 3097 3409 3106 3443
rect 2924 3392 3106 3409
rect 2664 3335 2850 3356
rect 2664 3301 2671 3335
rect 2671 3301 2839 3335
rect 2839 3301 2850 3335
rect 2664 3298 2850 3301
rect 2946 3066 3098 3122
<< metal2 >>
rect 2664 3690 2850 3692
rect 2664 3634 2684 3690
rect 2836 3634 2850 3690
rect 2664 3364 2850 3634
rect 2918 3446 3116 3454
rect 2918 3392 2924 3446
rect 3106 3392 3116 3446
rect 2656 3356 2860 3364
rect 2656 3298 2664 3356
rect 2850 3298 2860 3356
rect 2656 3290 2860 3298
rect 2918 3122 3116 3392
rect 2918 3066 2946 3122
rect 3098 3066 3116 3122
rect 2918 3060 3116 3066
<< labels >>
rlabel metal1 202 6635 301 6697 1 curgate
rlabel locali -880 7978 -840 8007 1 body
rlabel locali -240 3228 -160 3432 1 gnd1
rlabel locali -162 8062 -130 8134 1 gnd2
rlabel metal1 706 3206 938 3438 1 vp
rlabel locali 1368 1956 1458 2135 1 nwell
rlabel metal1 2994 3676 3044 3698 1 vout_p
rlabel metal1 2750 3042 2802 3066 1 vout_n
<< end >>
