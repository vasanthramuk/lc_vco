magic
tech sky130A
magscale 1 2
timestamp 1671515826
<< nwell >>
rect 1312 4027 3686 4314
rect 1312 1405 1683 4027
rect 3399 1405 3686 4027
rect 1312 1052 3686 1405
<< pwell >>
rect 276 8021 387 8079
rect 1683 1405 3399 4027
<< psubdiff >>
rect -326 505 -137 541
rect -326 403 -290 505
rect -183 403 -137 505
rect -326 368 -137 403
<< nsubdiff >>
rect 3499 4226 3641 4235
rect 1418 4204 3641 4226
rect 1418 4097 1445 4204
rect 3613 4131 3641 4204
rect 1420 1185 1445 4097
rect 1533 4097 3524 4131
rect 1533 1270 1555 4097
rect 3499 1270 3524 4097
rect 1533 1250 3524 1270
rect 3612 4094 3641 4131
rect 3612 1186 3634 4094
rect 3610 1185 3634 1186
rect 1420 1153 3634 1185
rect 3499 1151 3634 1153
<< psubdiffcont >>
rect -290 403 -183 505
<< nsubdiffcont >>
rect 1445 4131 3613 4204
rect 1445 1250 1533 4131
rect 3524 1250 3612 4131
rect 1445 1186 3612 1250
rect 1445 1185 3610 1186
<< polycont >>
rect 211 8013 276 8087
<< locali >>
rect 196 8087 300 8103
rect 196 8013 211 8087
rect 276 8079 300 8087
rect 276 8021 387 8079
rect 276 8013 300 8021
rect 196 7994 300 8013
rect 1420 4224 1549 4227
rect 1420 4204 3631 4224
rect 1420 1185 1445 4204
rect 3613 4131 3631 4204
rect 1533 4117 3524 4131
rect 1533 1265 1549 4117
rect 3502 1265 3524 4117
rect 1533 1250 3524 1265
rect 3612 1186 3631 4131
rect 3610 1185 3631 1186
rect 1420 1164 3631 1185
rect 1432 1160 3631 1164
rect 1432 1159 3626 1160
rect -312 505 -162 523
rect -312 403 -290 505
rect -183 403 -162 505
rect -312 381 -162 403
<< metal1 >>
rect 143 6515 341 6841
rect 143 6451 351 6515
use sky130_fd_pr__nfet_01v8_F8A7VK  sky130_fd_pr__nfet_01v8_F8A7VK_0
timestamp 1671513803
transform 1 0 243 0 1 3295
box -296 -3346 296 3346
use sky130_fd_pr__nfet_01v8_NFC7VK  sky130_fd_pr__nfet_01v8_NFC7VK_0
timestamp 1671513803
transform 1 0 241 0 1 8062
box -296 -1399 296 1399
use sky130_fd_pr__nfet_01v8_TPE47J  sky130_fd_pr__nfet_01v8_TPE47J_0
timestamp 1671515165
transform 1 0 2499 0 1 2712
box -683 -1119 683 1119
<< labels >>
rlabel psubdiffcont -282 406 -188 502 1 body
rlabel metal1 190 6615 312 6681 1 curgate
rlabel nsubdiffcont 1985 1185 2132 1241 1 nwell
rlabel space 102 7251 125 7329 1 GND!
rlabel space 102 5196 125 5262 1 GND!
rlabel space 360 5262 387 5314 1 vp
<< end >>
