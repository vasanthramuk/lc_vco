magic
tech sky130A
magscale 1 2
timestamp 1671528211
<< nwell >>
rect -1352 1268 1338 1534
rect -1352 -1268 -922 1268
rect 1004 -1268 1338 1268
rect -1352 -1546 1338 -1268
<< pwell >>
rect -922 -1268 1004 1268
<< nmos >>
rect -487 109 -287 909
rect -229 109 -29 909
rect 29 109 229 909
rect 287 109 487 909
rect -487 -909 -287 -109
rect -229 -909 -29 -109
rect 29 -909 229 -109
rect 287 -909 487 -109
<< ndiff >>
rect -545 897 -487 909
rect -545 121 -533 897
rect -499 121 -487 897
rect -545 109 -487 121
rect -287 897 -229 909
rect -287 121 -275 897
rect -241 121 -229 897
rect -287 109 -229 121
rect -29 897 29 909
rect -29 121 -17 897
rect 17 121 29 897
rect -29 109 29 121
rect 229 897 287 909
rect 229 121 241 897
rect 275 121 287 897
rect 229 109 287 121
rect 487 897 545 909
rect 487 121 499 897
rect 533 121 545 897
rect 487 109 545 121
rect -545 -121 -487 -109
rect -545 -897 -533 -121
rect -499 -897 -487 -121
rect -545 -909 -487 -897
rect -287 -121 -229 -109
rect -287 -897 -275 -121
rect -241 -897 -229 -121
rect -287 -909 -229 -897
rect -29 -121 29 -109
rect -29 -897 -17 -121
rect 17 -897 29 -121
rect -29 -909 29 -897
rect 229 -121 287 -109
rect 229 -897 241 -121
rect 275 -897 287 -121
rect 229 -909 287 -897
rect 487 -121 545 -109
rect 487 -897 499 -121
rect 533 -897 545 -121
rect 487 -909 545 -897
<< ndiffc >>
rect -533 121 -499 897
rect -275 121 -241 897
rect -17 121 17 897
rect 241 121 275 897
rect 499 121 533 897
rect -533 -897 -499 -121
rect -275 -897 -241 -121
rect -17 -897 17 -121
rect 241 -897 275 -121
rect 499 -897 533 -121
<< psubdiff >>
rect -647 1049 -551 1083
rect 551 1049 647 1083
rect -647 987 -613 1049
rect 613 987 647 1049
rect -647 -1049 -613 -987
rect 613 -1049 647 -987
rect -647 -1083 -551 -1049
rect 551 -1083 647 -1049
<< nsubdiff >>
rect 1096 1450 1264 1476
rect -1238 1434 1264 1450
rect -1238 1318 -1214 1434
rect 1202 1334 1264 1434
rect -1236 -1446 -1214 1318
rect -1090 1318 1118 1334
rect -1090 -1328 -1068 1318
rect 1094 -1328 1118 1318
rect -1090 -1348 1118 -1328
rect 1200 1322 1264 1334
rect 1200 -1348 1224 1322
rect 1202 -1446 1224 -1348
rect -1236 -1470 1224 -1446
<< psubdiffcont >>
rect -551 1049 551 1083
rect -647 -987 -613 987
rect 613 -987 647 987
rect -551 -1083 551 -1049
<< nsubdiffcont >>
rect -1214 1334 1202 1434
rect -1214 -1348 -1090 1334
rect 1118 -1348 1200 1334
rect -1214 -1446 1202 -1348
<< poly >>
rect -487 981 -287 997
rect -487 947 -471 981
rect -303 947 -287 981
rect -487 909 -287 947
rect -229 981 -29 997
rect -229 947 -213 981
rect -45 947 -29 981
rect -229 909 -29 947
rect 29 981 229 997
rect 29 947 45 981
rect 213 947 229 981
rect 29 909 229 947
rect 287 981 487 997
rect 287 947 303 981
rect 471 947 487 981
rect 287 909 487 947
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect -487 -947 -287 -909
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -487 -997 -287 -981
rect -229 -947 -29 -909
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect -229 -997 -29 -981
rect 29 -947 229 -909
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 29 -997 229 -981
rect 287 -947 487 -909
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 287 -997 487 -981
<< polycont >>
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
<< locali >>
rect -1254 1434 1238 1464
rect -1254 -1446 -1214 1434
rect 1202 1334 1238 1434
rect -1090 1330 1118 1334
rect -1090 -1306 -1004 1330
rect -647 1049 -551 1083
rect 551 1049 647 1083
rect -647 987 -613 1049
rect 613 987 647 1049
rect -487 947 -471 981
rect -303 947 -287 981
rect -229 947 -213 981
rect -45 947 -29 981
rect 29 947 45 981
rect 213 947 229 981
rect 287 947 303 981
rect 471 947 487 981
rect -533 897 -499 913
rect -275 897 -241 913
rect -533 105 -499 121
rect -17 897 17 913
rect 241 897 275 913
rect -275 105 -241 121
rect 499 897 533 913
rect -17 105 17 121
rect 241 105 275 121
rect 499 105 533 121
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect -533 -121 -499 -105
rect -275 -121 -241 -105
rect -17 -121 17 -105
rect -533 -913 -499 -897
rect 241 -121 275 -105
rect 499 -121 533 -105
rect -275 -913 -241 -897
rect -17 -913 17 -897
rect 241 -913 275 -897
rect 499 -913 533 -897
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 287 -981 303 -947
rect 471 -981 487 -947
rect -647 -1049 -613 -987
rect 613 -1049 647 -987
rect -647 -1083 -551 -1049
rect 551 -1083 647 -1049
rect 1080 -1306 1118 1330
rect -1090 -1348 1118 -1306
rect 1200 -1306 1238 1334
rect 1200 -1348 1240 -1306
rect 1202 -1446 1240 -1348
rect -1254 -1494 1240 -1446
rect -1254 -1498 -1004 -1494
<< viali >>
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect -534 746 -533 862
rect -533 746 -499 862
rect -499 746 -498 862
rect -18 744 -17 862
rect -17 744 17 862
rect 17 744 18 862
rect -274 266 -241 380
rect -241 266 -240 380
rect 498 744 499 862
rect 499 744 533 862
rect 533 744 534 862
rect 240 266 241 380
rect 241 266 274 380
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect -278 -378 -275 -262
rect -275 -378 -241 -262
rect -241 -378 -238 -262
rect -534 -868 -533 -752
rect -533 -868 -499 -752
rect -499 -868 -498 -752
rect 238 -374 241 -260
rect 241 -374 275 -260
rect 275 -374 278 -260
rect -18 -868 -17 -752
rect -17 -868 17 -752
rect 17 -868 18 -752
rect 498 -868 499 -752
rect 499 -868 533 -752
rect 533 -868 534 -752
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
<< metal1 >>
rect -483 981 -291 987
rect -483 947 -471 981
rect -303 947 -291 981
rect -483 941 -291 947
rect -225 981 -33 987
rect -225 947 -213 981
rect -45 947 -33 981
rect -225 941 -33 947
rect 33 981 225 987
rect 33 947 45 981
rect 213 947 225 981
rect 33 941 225 947
rect 291 981 483 987
rect 291 947 303 981
rect 471 947 483 981
rect 291 941 483 947
rect -546 862 548 874
rect -546 746 -534 862
rect -498 746 -18 862
rect -546 744 -18 746
rect 18 744 498 862
rect 534 744 548 862
rect -546 728 548 744
rect -290 380 294 390
rect -290 266 -274 380
rect -240 318 240 380
rect -240 266 -200 318
rect -290 262 -200 266
rect -48 266 240 318
rect 274 266 294 380
rect -48 262 294 266
rect -290 252 294 262
rect 34 77 226 78
rect -483 76 -291 77
rect -225 76 -33 77
rect 33 76 226 77
rect 291 76 483 77
rect -483 74 483 76
rect -483 71 40 74
rect 222 71 483 74
rect -483 37 -471 71
rect -303 37 -213 71
rect -45 37 40 71
rect 222 37 303 71
rect 471 37 483 71
rect -483 32 40 37
rect -483 31 -291 32
rect -225 31 -33 32
rect 33 31 40 32
rect 34 20 40 31
rect 222 32 483 37
rect 222 20 226 32
rect 291 31 483 32
rect 34 14 226 20
rect -226 -16 -28 -12
rect -483 -32 -291 -31
rect -226 -32 -220 -16
rect -483 -37 -220 -32
rect -34 -32 -28 -16
rect 33 -32 225 -31
rect 291 -32 483 -31
rect -34 -37 483 -32
rect -483 -71 -471 -37
rect -303 -71 -220 -37
rect -34 -71 45 -37
rect 213 -71 303 -37
rect 471 -71 483 -37
rect -483 -74 -220 -71
rect -34 -74 483 -71
rect -483 -77 -291 -74
rect -226 -76 -28 -74
rect -225 -77 -33 -76
rect 33 -77 225 -74
rect 291 -77 483 -74
rect -294 -250 300 -244
rect -294 -262 62 -250
rect -294 -378 -278 -262
rect -238 -306 62 -262
rect 214 -260 300 -250
rect 214 -306 238 -260
rect -238 -374 238 -306
rect 278 -374 300 -260
rect -238 -378 300 -374
rect -294 -390 300 -378
rect -544 -752 562 -740
rect -544 -868 -534 -752
rect -498 -868 -18 -752
rect 18 -868 498 -752
rect 534 -868 562 -752
rect -544 -890 562 -868
rect -483 -942 -291 -941
rect -225 -942 -33 -941
rect 33 -942 225 -941
rect 291 -942 483 -941
rect -483 -947 483 -942
rect -483 -981 -471 -947
rect -303 -981 -213 -947
rect -45 -981 45 -947
rect 213 -981 303 -947
rect 471 -981 483 -947
rect -483 -986 483 -981
rect -483 -987 -291 -986
rect -225 -987 -33 -986
rect 33 -987 225 -986
rect 291 -987 483 -986
<< via1 >>
rect -200 262 -48 318
rect 40 71 222 74
rect 40 37 45 71
rect 45 37 213 71
rect 213 37 222 71
rect 40 20 222 37
rect -220 -37 -34 -16
rect -220 -71 -213 -37
rect -213 -71 -45 -37
rect -45 -71 -34 -37
rect -220 -74 -34 -71
rect 62 -306 214 -250
<< metal2 >>
rect -220 318 -34 320
rect -220 262 -200 318
rect -48 262 -34 318
rect -220 -8 -34 262
rect 34 74 232 82
rect 34 20 40 74
rect 222 20 232 74
rect -228 -16 -24 -8
rect -228 -74 -220 -16
rect -34 -74 -24 -16
rect -228 -82 -24 -74
rect 34 -250 232 20
rect 34 -306 62 -250
rect 214 -306 232 -250
rect 34 -312 232 -306
<< properties >>
string FIXED_BBOX -630 -1066 630 1066
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 1 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
