* SPICE3 file created from trial.ext - technology: sky130A

X0 vp curgate curgate vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X1 vp curgate curgate vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X2 vp m3_5645_3434# m1_2766_4324# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3 vp m1_2766_4324# m3_5645_3434# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4 m3_5645_3434# m1_2766_4324# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5 vp m1_2766_4324# m3_5645_3434# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 m1_2766_4324# m3_5645_3434# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7 vp m3_5645_3434# m1_2766_4324# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8 m3_5645_3434# m1_2766_4324# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 m1_2766_4324# m3_5645_3434# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10 m1_2766_4324# vcntrl vp sky130_fd_pr__cap_var_lvt w=1e+07u l=500000u
X11 m3_5645_3434# vcntrl vp sky130_fd_pr__cap_var_lvt w=1e+07u l=500000u
X12 m4_n1090_3434# m1_2766_4324# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X13 m4_5645_3434# m3_5645_3434# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X14 m4_n1090_3434# m1_2766_4324# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X15 m4_5645_3434# m3_5645_3434# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X16 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X17 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X18 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X19 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X20 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
C0 m1_2766_4324# m4_n1090_3434# 88.15fF
C1 vcntrl m3_5645_3434# 2.52fF
C2 m3_5645_3434# m4_5645_3434# 88.14fF
C3 m3_5645_3434# m1_2766_4324# 5.64fF
C4 vcntrl m1_2766_4324# 2.50fF
C5 curgate vp 6.16fF **FLOATING
C6 m4_5645_3434# vp 4.01fF **FLOATING
C7 m4_n1090_3434# vp 4.02fF **FLOATING
C8 m1_2766_4324# vp 24.81fF **FLOATING
C9 vcntrl vp 9.09fF **FLOATING
C10 m3_5645_3434# vp 28.25fF **FLOATING
