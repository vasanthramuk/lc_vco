magic
tech sky130A
magscale 1 2
timestamp 1670838278
<< metal3 >>
rect -2413 2335 2412 2363
rect -2413 -2335 2328 2335
rect 2392 -2335 2412 2335
rect -2413 -2363 2412 -2335
<< via3 >>
rect 2328 -2335 2392 2335
<< mimcap >>
rect -2313 2223 2213 2263
rect -2313 -2223 -2273 2223
rect 2173 -2223 2213 2223
rect -2313 -2263 2213 -2223
<< mimcapcontact >>
rect -2273 -2223 2173 2223
<< metal4 >>
rect 2312 2335 2408 2351
rect -2274 2223 2174 2224
rect -2274 -2223 -2273 2223
rect 2173 -2223 2174 2223
rect -2274 -2224 2174 -2223
rect 2312 -2335 2328 2335
rect 2392 -2335 2408 2335
rect 2312 -2351 2408 -2335
<< properties >>
string FIXED_BBOX -2413 -2363 2313 2363
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 22.63 l 22.63 val 1.041k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
