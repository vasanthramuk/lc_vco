magic
tech sky130A
magscale 1 2
timestamp 1671439731
<< locali >>
rect 3054 2182 3424 2190
rect 3054 2136 3174 2182
rect 3166 2126 3174 2136
rect 3292 2136 3424 2182
rect 3292 2126 3300 2136
rect 3166 2118 3300 2126
rect -1698 -92 -1570 102
rect -306 -16 18 54
rect 3228 -2 3428 130
rect 3138 -40 3428 -2
rect 3138 -104 3188 -40
rect 3282 -104 3428 -40
rect 3138 -158 3428 -104
<< viali >>
rect 3174 2126 3292 2182
rect 2424 2006 2592 2058
rect 3912 758 4078 810
rect 3188 -104 3282 -40
<< metal1 >>
rect 2705 2336 3765 4251
rect 2412 2058 2610 2074
rect 2412 2006 2424 2058
rect 2592 2006 2610 2058
rect 2412 2000 2610 2006
rect 2412 1948 2608 2000
rect 2740 1628 2990 2268
rect 3160 2190 3308 2196
rect 3160 2120 3168 2190
rect 3302 2120 3308 2190
rect 3160 2112 3308 2120
rect 3490 1628 3740 2268
rect 2466 841 2518 862
rect 3953 852 4087 911
rect 2425 798 2559 841
rect 3890 810 4087 852
rect 2412 733 2652 798
rect 3890 758 3912 810
rect 4078 758 4087 810
rect 3890 733 4087 758
rect 2412 656 4087 733
rect 2421 487 4087 656
rect 2421 457 3715 487
rect 2923 355 3715 457
rect 3059 353 3715 355
rect 3127 347 3715 353
rect -406 160 118 324
rect 3174 -40 3298 -30
rect 3174 -104 3188 -40
rect 3282 -104 3298 -40
rect 3174 -118 3298 -104
<< via1 >>
rect 3168 2182 3302 2190
rect 3168 2126 3174 2182
rect 3174 2126 3292 2182
rect 3292 2126 3302 2182
rect 3168 2120 3302 2126
rect 3188 -104 3282 -40
<< metal2 >>
rect 2622 5286 2990 5524
rect 2622 4986 2686 5286
rect 2922 4986 2990 5286
rect 2622 4196 2990 4986
rect 3462 5286 3830 5524
rect 3462 4986 3532 5286
rect 3768 4986 3830 5286
rect 3462 4196 3830 4986
rect 3158 2190 3312 2200
rect 3158 2120 3168 2190
rect 3302 2120 3312 2190
rect 3158 2110 3312 2120
rect 3174 -40 3296 -30
rect 3174 -104 3188 -40
rect 3282 -104 3296 -40
rect 3174 -118 3296 -104
<< via2 >>
rect 2686 4986 2922 5286
rect 3532 4986 3768 5286
rect 3170 2122 3296 2188
rect 3188 -104 3282 -40
<< metal3 >>
rect 1972 5286 2990 5572
rect 1972 4986 2686 5286
rect 2922 4986 2990 5286
rect 1972 4778 2990 4986
rect 3462 5286 4500 5572
rect 3462 4986 3532 5286
rect 3768 4986 4500 5286
rect 3462 4776 4500 4986
rect -1074 3450 863 4201
rect 5645 3434 7605 4201
rect 3158 2188 3312 2200
rect 3158 2122 3170 2188
rect 3296 2122 3312 2188
rect 3158 2110 3312 2122
rect 3170 -40 3294 2110
rect 3170 -104 3188 -40
rect 3282 -104 3294 -40
rect 3170 -130 3294 -104
<< metal4 >>
rect -1090 4200 870 4201
rect 5645 4200 7605 4201
rect -1090 3446 7605 4200
rect -1090 3434 870 3446
rect 5645 3434 7605 3446
use sky130_fd_pr__cap_mim_m3_1_8UNQ5L  sky130_fd_pr__cap_mim_m3_1_8UNQ5L_0
timestamp 1670838128
transform 1 0 30 0 1 1477
box -2413 -2363 2412 2363
use sky130_fd_pr__cap_mim_m3_1_8UNQ5L  sky130_fd_pr__cap_mim_m3_1_8UNQ5L_1
timestamp 1670838128
transform -1 0 6392 0 -1 1477
box -2413 -2363 2412 2363
use sky130_fd_pr__cap_mim_m3_1_8UNQ5L  sky130_fd_pr__cap_mim_m3_1_8UNQ5L_2
timestamp 1670838128
transform 1 0 30 0 1 6289
box -2413 -2363 2412 2363
use sky130_fd_pr__cap_mim_m3_1_8UNQ5L  sky130_fd_pr__cap_mim_m3_1_8UNQ5L_3
timestamp 1670838128
transform -1 0 6392 0 -1 6289
box -2413 -2363 2412 2363
use sky130_fd_pr__cap_var_lvt_E5Z3X6  sky130_fd_pr__cap_var_lvt_E5Z3X6_0
timestamp 1671439258
transform 1 0 2812 0 1 3292
box -293 -1201 293 1201
use sky130_fd_pr__cap_var_lvt_E5Z3X6  sky130_fd_pr__cap_var_lvt_E5Z3X6_1
timestamp 1671439258
transform 1 0 3655 0 1 3292
box -293 -1201 293 1201
use sky130_fd_pr__nfet_01v8_F8A7VK  sky130_fd_pr__nfet_01v8_F8A7VK_0
timestamp 1671089082
transform 0 1 3293 -1 0 243
box -296 -3571 371 3346
use sky130_fd_pr__nfet_01v8_NFC7VK  sky130_fd_pr__nfet_01v8_NFC7VK_0
timestamp 1671430078
transform 0 1 -1636 -1 0 243
box -449 -1399 331 1399
use sky130_fd_pr__nfet_01v8_TPE47J  sky130_fd_pr__nfet_01v8_TPE47J_0
timestamp 1671089082
transform 0 1 3254 -1 0 1404
box -683 -1119 683 1119
use sky130_fd_pr__nfet_01v8_VYRQW9  sky130_fd_pr__nfet_01v8_VYRQW9_0
timestamp 1670822484
transform 0 1 3220 -1 0 1149
box 0 0 1 1
<< labels >>
rlabel metal1 3140 530 3532 694 1 vp
rlabel metal1 -258 192 -48 310 1 curgate
rlabel space 2979 1511 3133 1562 1 vout_m
rlabel space 3346 1268 3528 1319 1 vout_p
rlabel locali -1646 -72 -1620 -36 1 gnd
port 1 n
rlabel locali 3304 -124 3334 -70 1 gnd
rlabel metal1 3112 2888 3368 3624 1 vcntrl
rlabel metal4 3024 3762 3452 3998 1 VDD
<< end >>
