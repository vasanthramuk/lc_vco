magic
tech sky130A
magscale 1 2
timestamp 1670046323
<< error_p >>
rect -70 6500 -10 10700
rect 10 6500 70 10700
rect -70 2200 -10 6400
rect 10 2200 70 6400
rect -70 -2100 -10 2100
rect 10 -2100 70 2100
rect -70 -6400 -10 -2200
rect 10 -6400 70 -2200
rect -70 -10700 -10 -6500
rect 10 -10700 70 -6500
<< metal3 >>
rect -6309 10672 -10 10700
rect -6309 6528 -94 10672
rect -30 6528 -10 10672
rect -6309 6500 -10 6528
rect 10 10672 6309 10700
rect 10 6528 6225 10672
rect 6289 6528 6309 10672
rect 10 6500 6309 6528
rect -6309 6372 -10 6400
rect -6309 2228 -94 6372
rect -30 2228 -10 6372
rect -6309 2200 -10 2228
rect 10 6372 6309 6400
rect 10 2228 6225 6372
rect 6289 2228 6309 6372
rect 10 2200 6309 2228
rect -6309 2072 -10 2100
rect -6309 -2072 -94 2072
rect -30 -2072 -10 2072
rect -6309 -2100 -10 -2072
rect 10 2072 6309 2100
rect 10 -2072 6225 2072
rect 6289 -2072 6309 2072
rect 10 -2100 6309 -2072
rect -6309 -2228 -10 -2200
rect -6309 -6372 -94 -2228
rect -30 -6372 -10 -2228
rect -6309 -6400 -10 -6372
rect 10 -2228 6309 -2200
rect 10 -6372 6225 -2228
rect 6289 -6372 6309 -2228
rect 10 -6400 6309 -6372
rect -6309 -6528 -10 -6500
rect -6309 -10672 -94 -6528
rect -30 -10672 -10 -6528
rect -6309 -10700 -10 -10672
rect 10 -6528 6309 -6500
rect 10 -10672 6225 -6528
rect 6289 -10672 6309 -6528
rect 10 -10700 6309 -10672
<< via3 >>
rect -94 6528 -30 10672
rect 6225 6528 6289 10672
rect -94 2228 -30 6372
rect 6225 2228 6289 6372
rect -94 -2072 -30 2072
rect 6225 -2072 6289 2072
rect -94 -6372 -30 -2228
rect 6225 -6372 6289 -2228
rect -94 -10672 -30 -6528
rect 6225 -10672 6289 -6528
<< mimcap >>
rect -6209 10560 -209 10600
rect -6209 6640 -6169 10560
rect -249 6640 -209 10560
rect -6209 6600 -209 6640
rect 110 10560 6110 10600
rect 110 6640 150 10560
rect 6070 6640 6110 10560
rect 110 6600 6110 6640
rect -6209 6260 -209 6300
rect -6209 2340 -6169 6260
rect -249 2340 -209 6260
rect -6209 2300 -209 2340
rect 110 6260 6110 6300
rect 110 2340 150 6260
rect 6070 2340 6110 6260
rect 110 2300 6110 2340
rect -6209 1960 -209 2000
rect -6209 -1960 -6169 1960
rect -249 -1960 -209 1960
rect -6209 -2000 -209 -1960
rect 110 1960 6110 2000
rect 110 -1960 150 1960
rect 6070 -1960 6110 1960
rect 110 -2000 6110 -1960
rect -6209 -2340 -209 -2300
rect -6209 -6260 -6169 -2340
rect -249 -6260 -209 -2340
rect -6209 -6300 -209 -6260
rect 110 -2340 6110 -2300
rect 110 -6260 150 -2340
rect 6070 -6260 6110 -2340
rect 110 -6300 6110 -6260
rect -6209 -6640 -209 -6600
rect -6209 -10560 -6169 -6640
rect -249 -10560 -209 -6640
rect -6209 -10600 -209 -10560
rect 110 -6640 6110 -6600
rect 110 -10560 150 -6640
rect 6070 -10560 6110 -6640
rect 110 -10600 6110 -10560
<< mimcapcontact >>
rect -6169 6640 -249 10560
rect 150 6640 6070 10560
rect -6169 2340 -249 6260
rect 150 2340 6070 6260
rect -6169 -1960 -249 1960
rect 150 -1960 6070 1960
rect -6169 -6260 -249 -2340
rect 150 -6260 6070 -2340
rect -6169 -10560 -249 -6640
rect 150 -10560 6070 -6640
<< metal4 >>
rect -3261 10561 -3157 10750
rect -141 10688 -37 10750
rect -141 10672 -14 10688
rect -6170 10560 -248 10561
rect -6170 6640 -6169 10560
rect -249 6640 -248 10560
rect -6170 6639 -248 6640
rect -3261 6261 -3157 6639
rect -141 6528 -94 10672
rect -30 6528 -14 10672
rect 3058 10561 3162 10750
rect 6178 10688 6282 10750
rect 6178 10672 6305 10688
rect 149 10560 6071 10561
rect 149 6640 150 10560
rect 6070 6640 6071 10560
rect 149 6639 6071 6640
rect -141 6512 -14 6528
rect -141 6388 -37 6512
rect -141 6372 -14 6388
rect -6170 6260 -248 6261
rect -6170 2340 -6169 6260
rect -249 2340 -248 6260
rect -6170 2339 -248 2340
rect -3261 1961 -3157 2339
rect -141 2228 -94 6372
rect -30 2228 -14 6372
rect 3058 6261 3162 6639
rect 6178 6528 6225 10672
rect 6289 6528 6305 10672
rect 6178 6512 6305 6528
rect 6178 6388 6282 6512
rect 6178 6372 6305 6388
rect 149 6260 6071 6261
rect 149 2340 150 6260
rect 6070 2340 6071 6260
rect 149 2339 6071 2340
rect -141 2212 -14 2228
rect -141 2088 -37 2212
rect -141 2072 -14 2088
rect -6170 1960 -248 1961
rect -6170 -1960 -6169 1960
rect -249 -1960 -248 1960
rect -6170 -1961 -248 -1960
rect -3261 -2339 -3157 -1961
rect -141 -2072 -94 2072
rect -30 -2072 -14 2072
rect 3058 1961 3162 2339
rect 6178 2228 6225 6372
rect 6289 2228 6305 6372
rect 6178 2212 6305 2228
rect 6178 2088 6282 2212
rect 6178 2072 6305 2088
rect 149 1960 6071 1961
rect 149 -1960 150 1960
rect 6070 -1960 6071 1960
rect 149 -1961 6071 -1960
rect -141 -2088 -14 -2072
rect -141 -2212 -37 -2088
rect -141 -2228 -14 -2212
rect -6170 -2340 -248 -2339
rect -6170 -6260 -6169 -2340
rect -249 -6260 -248 -2340
rect -6170 -6261 -248 -6260
rect -3261 -6639 -3157 -6261
rect -141 -6372 -94 -2228
rect -30 -6372 -14 -2228
rect 3058 -2339 3162 -1961
rect 6178 -2072 6225 2072
rect 6289 -2072 6305 2072
rect 6178 -2088 6305 -2072
rect 6178 -2212 6282 -2088
rect 6178 -2228 6305 -2212
rect 149 -2340 6071 -2339
rect 149 -6260 150 -2340
rect 6070 -6260 6071 -2340
rect 149 -6261 6071 -6260
rect -141 -6388 -14 -6372
rect -141 -6512 -37 -6388
rect -141 -6528 -14 -6512
rect -6170 -6640 -248 -6639
rect -6170 -10560 -6169 -6640
rect -249 -10560 -248 -6640
rect -6170 -10561 -248 -10560
rect -3261 -10750 -3157 -10561
rect -141 -10672 -94 -6528
rect -30 -10672 -14 -6528
rect 3058 -6639 3162 -6261
rect 6178 -6372 6225 -2228
rect 6289 -6372 6305 -2228
rect 6178 -6388 6305 -6372
rect 6178 -6512 6282 -6388
rect 6178 -6528 6305 -6512
rect 149 -6640 6071 -6639
rect 149 -10560 150 -6640
rect 6070 -10560 6071 -6640
rect 149 -10561 6071 -10560
rect -141 -10688 -14 -10672
rect -141 -10750 -37 -10688
rect 3058 -10750 3162 -10561
rect 6178 -10672 6225 -6528
rect 6289 -10672 6305 -6528
rect 6178 -10688 6305 -10672
rect 6178 -10750 6282 -10688
<< properties >>
string FIXED_BBOX 10 6500 6210 10700
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 20 val 1.219k carea 2.00 cperi 0.19 nx 2 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
