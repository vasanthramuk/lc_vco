magic
tech sky130A
magscale 1 2
timestamp 1670824296
<< pwell >>
rect -683 -610 683 610
<< nmos >>
rect -487 -400 -287 400
rect -229 -400 -29 400
rect 29 -400 229 400
rect 287 -400 487 400
<< ndiff >>
rect -545 388 -487 400
rect -545 -388 -533 388
rect -499 -388 -487 388
rect -545 -400 -487 -388
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
rect 487 388 545 400
rect 487 -388 499 388
rect 533 -388 545 388
rect 487 -400 545 -388
<< ndiffc >>
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
<< psubdiff >>
rect -647 540 -551 574
rect 551 540 647 574
rect -647 478 -613 540
rect 613 478 647 540
rect -647 -540 -613 -478
rect 613 -540 647 -478
rect -647 -574 -551 -540
rect 551 -574 647 -540
<< psubdiffcont >>
rect -551 540 551 574
rect -647 -478 -613 478
rect 613 -478 647 478
rect -551 -574 551 -540
<< poly >>
rect -487 472 -287 488
rect -487 438 -471 472
rect -303 438 -287 472
rect -487 400 -287 438
rect -229 472 -29 488
rect -229 438 -213 472
rect -45 438 -29 472
rect -229 400 -29 438
rect 29 472 229 488
rect 29 438 45 472
rect 213 438 229 472
rect 29 400 229 438
rect 287 472 487 488
rect 287 438 303 472
rect 471 438 487 472
rect 287 400 487 438
rect -487 -438 -287 -400
rect -487 -472 -471 -438
rect -303 -472 -287 -438
rect -487 -488 -287 -472
rect -229 -438 -29 -400
rect -229 -472 -213 -438
rect -45 -472 -29 -438
rect -229 -488 -29 -472
rect 29 -438 229 -400
rect 29 -472 45 -438
rect 213 -472 229 -438
rect 29 -488 229 -472
rect 287 -438 487 -400
rect 287 -472 303 -438
rect 471 -472 487 -438
rect 287 -488 487 -472
<< polycont >>
rect -471 438 -303 472
rect -213 438 -45 472
rect 45 438 213 472
rect 303 438 471 472
rect -471 -472 -303 -438
rect -213 -472 -45 -438
rect 45 -472 213 -438
rect 303 -472 471 -438
<< locali >>
rect -647 540 -551 574
rect 551 540 647 574
rect -647 478 -613 540
rect 613 478 647 540
rect -487 438 -471 472
rect -303 438 -287 472
rect -229 438 -213 472
rect -45 438 -29 472
rect 29 438 45 472
rect 213 438 229 472
rect 287 438 303 472
rect 471 438 487 472
rect -533 388 -499 404
rect -533 -404 -499 -388
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
rect 499 388 533 404
rect 499 -404 533 -388
rect -487 -472 -471 -438
rect -303 -472 -287 -438
rect -229 -472 -213 -438
rect -45 -472 -29 -438
rect 29 -472 45 -438
rect 213 -472 229 -438
rect 287 -472 303 -438
rect 471 -472 487 -438
rect -647 -540 -613 -478
rect 613 -540 647 -478
rect -647 -574 -551 -540
rect 551 -574 647 -540
<< viali >>
rect -471 438 -303 472
rect -213 438 -45 472
rect 45 438 213 472
rect 303 438 471 472
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect -471 -472 -303 -438
rect -213 -472 -45 -438
rect 45 -472 213 -438
rect 303 -472 471 -438
<< metal1 >>
rect -483 472 -291 478
rect -483 438 -471 472
rect -303 438 -291 472
rect -483 432 -291 438
rect -225 472 -33 478
rect -225 438 -213 472
rect -45 438 -33 472
rect -225 432 -33 438
rect 33 472 225 478
rect 33 438 45 472
rect 213 438 225 472
rect 33 432 225 438
rect 291 472 483 478
rect 291 438 303 472
rect 471 438 483 472
rect 291 432 483 438
rect -539 388 -493 400
rect -539 -388 -533 388
rect -499 -388 -493 388
rect -539 -400 -493 -388
rect -281 388 -235 400
rect -281 -388 -275 388
rect -241 -388 -235 388
rect -281 -400 -235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 235 388 281 400
rect 235 -388 241 388
rect 275 -388 281 388
rect 235 -400 281 -388
rect 493 388 539 400
rect 493 -388 499 388
rect 533 -388 539 388
rect 493 -400 539 -388
rect -483 -438 -291 -432
rect -483 -472 -471 -438
rect -303 -472 -291 -438
rect -483 -478 -291 -472
rect -225 -438 -33 -432
rect -225 -472 -213 -438
rect -45 -472 -33 -438
rect -225 -478 -33 -472
rect 33 -438 225 -432
rect 33 -472 45 -438
rect 213 -472 225 -438
rect 33 -478 225 -472
rect 291 -438 483 -432
rect 291 -472 303 -438
rect 471 -472 483 -438
rect 291 -478 483 -472
<< properties >>
string FIXED_BBOX -630 -557 630 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
