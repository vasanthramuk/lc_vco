magic
tech sky130A
magscale 1 2
timestamp 1671533087
<< psubdiff >>
rect -919 8014 -802 8039
rect -919 7967 -887 8014
rect -829 7967 -802 8014
rect -919 7943 -802 7967
<< psubdiffcont >>
rect -887 7967 -829 8014
<< locali >>
rect -910 8014 -807 8037
rect -910 7967 -887 8014
rect -829 7967 -807 8014
rect -218 7988 52 8214
rect -910 7948 -807 7967
rect 2230 4234 2282 4240
rect 2230 4118 2236 4234
rect 2272 4118 2282 4234
rect 2230 4112 2282 4118
rect 3490 4236 3540 4240
rect 3490 4118 3496 4236
rect 3532 4118 3540 4236
rect 3490 4112 3540 4118
rect -370 2768 50 3820
rect 2228 2620 2282 2626
rect 2228 2504 2236 2620
rect 2272 2504 2282 2620
rect 2228 2496 2282 2504
rect 3487 2619 3539 2622
rect 3487 2503 3496 2619
rect 3532 2503 3539 2619
rect 3487 2495 3539 2503
rect 1311 1901 1880 2190
<< viali >>
rect 2236 4118 2272 4234
rect 3496 4118 3532 4236
rect 2236 2504 2272 2620
rect 3496 2503 3532 2619
<< metal1 >>
rect 146 6462 337 6876
rect 1200 4234 2427 4248
rect 1200 4118 2236 4234
rect 2272 4118 2427 4234
rect 1200 4099 2427 4118
rect 3402 4236 3548 4246
rect 3402 4118 3496 4236
rect 3532 4118 3548 4236
rect 3402 4100 3548 4118
rect 582 3836 930 3840
rect 1200 3836 1474 4099
rect 368 2750 1479 3836
rect 2934 3640 3086 3724
rect 2716 3016 2844 3086
rect 872 2749 1479 2750
rect 1198 2630 1479 2749
rect 3399 2630 3530 2631
rect 1198 2620 2432 2630
rect 1198 2504 2236 2620
rect 2272 2504 2432 2620
rect 1198 2482 2432 2504
rect 3399 2619 3548 2630
rect 3399 2503 3496 2619
rect 3532 2503 3548 2619
rect 3399 2481 3548 2503
rect 3480 2480 3548 2481
use sky130_fd_pr__nfet_01v8_F8A7VK  sky130_fd_pr__nfet_01v8_F8A7VK_0
timestamp 1671525571
transform 1 0 243 0 1 3293
box -296 -3346 296 3346
use sky130_fd_pr__nfet_01v8_NFC7VK  sky130_fd_pr__nfet_01v8_NFC7VK_0
timestamp 1671525571
transform 1 0 241 0 1 8098
box -296 -1399 296 1399
use sky130_fd_pr__nfet_01v8_TPE47J  sky130_fd_pr__nfet_01v8_TPE47J_0
timestamp 1671528211
transform 1 0 2884 0 1 3372
box -1352 -1546 1338 1534
<< labels >>
rlabel metal1 202 6635 301 6697 1 curgate
rlabel locali -880 7978 -840 8007 1 body
rlabel metal1 2750 3042 2802 3066 1 vout_n
rlabel metal1 2994 3676 3044 3698 1 vout_p
rlabel locali 1368 1956 1458 2135 1 nwell
rlabel locali -240 3228 -160 3432 1 gnd1
rlabel locali -162 8062 -130 8134 1 gnd2
rlabel metal1 706 3206 938 3438 1 vp
<< end >>
