* SPICE3 file created from sonamutha.ext - technology: sky130A

X0 vp curgate curgate vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X1 vp curgate curgate vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X2 vp m3_5645_4434# m3_5645_4434# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3 vp m3_5645_4434# m3_5645_4434# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4 m3_5645_4434# m3_5645_4434# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5 vp m3_5645_4434# m3_5645_4434# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 m3_5645_4434# m3_5645_4434# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7 vp m3_5645_4434# m3_5645_4434# vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8 m3_5645_4434# m3_5645_4434# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 m3_5645_4434# m3_5645_4434# vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10 m3_5645_4434# m1_2705_3336# vp sky130_fd_pr__cap_var_lvt w=1e+07u l=500000u
X11 m3_5645_4434# m1_2705_3336# vp sky130_fd_pr__cap_var_lvt w=1e+07u l=500000u
X12 m3_5645_4434# m3_5645_4434# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X13 m3_5645_4434# m3_5645_4434# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X14 m3_5645_4434# m3_5645_4434# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X15 m3_5645_4434# m3_5645_4434# sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X16 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X17 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X18 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X19 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X20 vp curgate vp vp sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
C0 m1_2705_3336# m3_5645_4434# 5.33fF
C1 curgate vp 6.22fF **FLOATING
C2 m3_5645_4434# vp 63.81fF **FLOATING
C3 m1_2705_3336# vp 9.14fF **FLOATING
C4 sky130_fd_pr__nfet_01v8_TPE47J_0/w_n1018_n1448# vp 7.16fF **FLOATING
