* SPICE3 file created from inductor.ext - technology: sky130A

C0 sky130_fd_pr__rf_test_coil1_0/m2_n4123_n14504# VSUBS 206.22fF **FLOATING
