magic
tech sky130A
magscale 1 2
timestamp 1671513803
<< error_p >>
rect -84 -1233 84 -1227
rect -84 -1255 -78 -1233
rect 78 -1255 84 -1233
rect -84 -1261 84 -1255
<< pwell >>
rect -296 -1399 296 1399
<< nmos >>
rect -100 109 100 1189
rect -100 -1189 100 -109
<< ndiff >>
rect -158 1177 -100 1189
rect -158 121 -146 1177
rect -112 121 -100 1177
rect -158 109 -100 121
rect 100 1177 158 1189
rect 100 121 112 1177
rect 146 121 158 1177
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -1177 -146 -121
rect -112 -1177 -100 -121
rect -158 -1189 -100 -1177
rect 100 -121 158 -109
rect 100 -1177 112 -121
rect 146 -1177 158 -121
rect 100 -1189 158 -1177
<< ndiffc >>
rect -146 121 -112 1177
rect 112 121 146 1177
rect -146 -1177 -112 -121
rect 112 -1177 146 -121
<< psubdiff >>
rect -260 1329 -164 1363
rect 164 1329 260 1363
rect -260 1267 -226 1329
rect 226 1267 260 1329
rect -260 -1329 -226 -1267
rect 226 -1329 260 -1267
rect -260 -1363 -164 -1329
rect 164 -1363 260 -1329
<< psubdiffcont >>
rect -164 1329 164 1363
rect -260 -1267 -226 1267
rect 226 -1267 260 1267
rect -164 -1363 164 -1329
<< poly >>
rect -100 1261 100 1277
rect -100 1227 -84 1261
rect 84 1227 100 1261
rect -100 1189 100 1227
rect -100 -109 100 109
rect -100 -1227 100 -1189
rect -100 -1261 -84 -1227
rect 84 -1261 100 -1227
rect -100 -1277 100 -1261
<< polycont >>
rect -84 1227 84 1261
rect -84 -1261 84 -1227
<< locali >>
rect -260 1329 -164 1363
rect 164 1329 260 1363
rect -260 1267 -226 1329
rect 226 1267 260 1329
rect -100 1227 -84 1261
rect 84 1227 100 1261
rect -146 1177 -112 1193
rect -146 -121 -112 121
rect -146 -1193 -112 -1177
rect 112 1177 146 1193
rect 112 -121 146 121
rect 112 -1193 146 -1177
rect -100 -1261 -84 -1227
rect 84 -1261 100 -1227
rect -260 -1329 -226 -1267
rect 226 -1329 260 -1267
rect -260 -1363 -164 -1329
rect 164 -1363 260 -1329
<< viali >>
rect -84 -1261 84 -1227
<< properties >>
string FIXED_BBOX -243 -1346 243 1346
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.4 l 1 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
