magic
tech sky130A
magscale 1 2
timestamp 1671445945
<< locali >>
rect 3054 3182 3424 3190
rect 3054 3136 3174 3182
rect 3166 3126 3174 3136
rect 3292 3136 3424 3182
rect 3292 3126 3300 3136
rect 3166 3118 3300 3126
rect -1698 -92 -1570 102
rect -306 -16 18 54
rect 3228 -2 3428 130
rect 3138 -40 3428 -2
rect 3138 -104 3188 -40
rect 3282 -104 3428 -40
rect 3138 -158 3428 -104
<< viali >>
rect 3174 3126 3292 3182
rect 3188 -104 3282 -40
<< metal1 >>
rect 2705 3336 3765 5251
rect 2740 2628 2990 3268
rect 3160 3190 3308 3196
rect 3160 3120 3168 3190
rect 3302 3120 3308 3190
rect 3160 3112 3308 3120
rect 3490 2628 3740 3268
rect 2867 2590 2946 2628
rect 2868 2500 2946 2590
rect 2867 2019 2946 2500
rect 3552 2018 3620 2628
rect 3953 1246 4087 1260
rect 2412 1152 2600 1178
rect 2412 798 2608 1152
rect 3892 852 4087 1246
rect 2412 733 2652 798
rect 3890 733 4087 852
rect 2412 656 4087 733
rect 2421 487 4087 656
rect 2421 457 3715 487
rect 2923 355 3715 457
rect 3059 353 3715 355
rect 3127 347 3715 353
rect -406 160 118 324
rect 3174 -40 3298 -30
rect 3174 -104 3188 -40
rect 3282 -104 3298 -40
rect 3174 -118 3298 -104
<< via1 >>
rect 3168 3182 3302 3190
rect 3168 3126 3174 3182
rect 3174 3126 3292 3182
rect 3292 3126 3302 3182
rect 3168 3120 3302 3126
rect 3188 -104 3282 -40
<< metal2 >>
rect 2622 6286 2990 6524
rect 2622 5986 2686 6286
rect 2922 5986 2990 6286
rect 2622 5196 2990 5986
rect 3462 6286 3830 6524
rect 3462 5986 3532 6286
rect 3768 5986 3830 6286
rect 3462 5196 3830 5986
rect 3158 3190 3312 3200
rect 3158 3120 3168 3190
rect 3302 3120 3312 3190
rect 3158 3110 3312 3120
rect 3174 -40 3296 -30
rect 3174 -104 3188 -40
rect 3282 -104 3296 -40
rect 3174 -118 3296 -104
<< via2 >>
rect 2686 5986 2922 6286
rect 3532 5986 3768 6286
rect 3170 3122 3296 3188
rect 3188 -104 3282 -40
<< metal3 >>
rect 1972 6286 2990 6572
rect 1972 5986 2686 6286
rect 2922 5986 2990 6286
rect 1972 5778 2990 5986
rect 3462 6286 4500 6572
rect 3462 5986 3532 6286
rect 3768 5986 4500 6286
rect 3462 5776 4500 5986
rect -1074 4450 863 5201
rect 5645 4434 7605 5201
rect 3158 3188 3312 3200
rect 3158 3122 3170 3188
rect 3296 3122 3312 3188
rect 3158 3110 3312 3122
rect 3170 -40 3294 3110
rect 3170 -104 3188 -40
rect 3282 -104 3294 -40
rect 3170 -130 3294 -104
<< metal4 >>
rect -1090 5200 870 5201
rect 5645 5200 7605 5201
rect -1072 4446 842 5200
rect -1090 4434 870 4446
rect -1072 4426 842 4434
rect 5636 4430 7608 5200
use sky130_fd_pr__cap_mim_m3_1_8UNQ5L  sky130_fd_pr__cap_mim_m3_1_8UNQ5L_0
timestamp 1670838128
transform 1 0 30 0 1 2477
box -2413 -2363 2412 2363
use sky130_fd_pr__cap_mim_m3_1_8UNQ5L  sky130_fd_pr__cap_mim_m3_1_8UNQ5L_1
timestamp 1670838128
transform -1 0 6392 0 -1 2477
box -2413 -2363 2412 2363
use sky130_fd_pr__cap_mim_m3_1_8UNQ5L  sky130_fd_pr__cap_mim_m3_1_8UNQ5L_2
timestamp 1670838128
transform 1 0 30 0 1 7289
box -2413 -2363 2412 2363
use sky130_fd_pr__cap_mim_m3_1_8UNQ5L  sky130_fd_pr__cap_mim_m3_1_8UNQ5L_3
timestamp 1670838128
transform -1 0 6392 0 -1 7289
box -2413 -2363 2412 2363
use sky130_fd_pr__cap_var_lvt_E5Z3X6  sky130_fd_pr__cap_var_lvt_E5Z3X6_0
timestamp 1671439258
transform 1 0 2812 0 1 4292
box -293 -1201 293 1201
use sky130_fd_pr__cap_var_lvt_E5Z3X6  sky130_fd_pr__cap_var_lvt_E5Z3X6_1
timestamp 1671439258
transform 1 0 3655 0 1 4292
box -293 -1201 293 1201
use sky130_fd_pr__nfet_01v8_F8A7VK  sky130_fd_pr__nfet_01v8_F8A7VK_0
timestamp 1671089082
transform 0 1 3293 -1 0 243
box -296 -3571 371 3346
use sky130_fd_pr__nfet_01v8_NFC7VK  sky130_fd_pr__nfet_01v8_NFC7VK_0
timestamp 1671430078
transform 0 1 -1636 -1 0 243
box -449 -1399 331 1399
use sky130_fd_pr__nfet_01v8_TPE47J  sky130_fd_pr__nfet_01v8_TPE47J_0
timestamp 1671443024
transform 0 1 3254 -1 0 1804
box -1018 -1448 890 1388
use sky130_fd_pr__nfet_01v8_VYRQW9  sky130_fd_pr__nfet_01v8_VYRQW9_0
timestamp 1670822484
transform 0 1 3220 -1 0 1149
box 0 0 1 1
<< labels >>
rlabel metal1 3406 560 3653 669 1 vp
rlabel locali 3316 -119 3398 -62 1 gnd
rlabel metal1 -204 173 -87 202 1 curgate
rlabel space 2978 1904 3114 1958 1 vout_m
rlabel space 3378 1670 3498 1718 1 vout_n
rlabel metal4 -370 4804 32 4994 1 VDD!
rlabel metal4 6408 4804 7170 5010 1 VDD!
<< end >>
