magic
tech sky130A
magscale 1 2
timestamp 1670733274
<< pwell >>
rect -396 -1399 396 1399
<< nmos >>
rect -200 109 200 1189
rect -200 -1189 200 -109
<< ndiff >>
rect -258 1177 -200 1189
rect -258 121 -246 1177
rect -212 121 -200 1177
rect -258 109 -200 121
rect 200 1177 258 1189
rect 200 121 212 1177
rect 246 121 258 1177
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -1177 -246 -121
rect -212 -1177 -200 -121
rect -258 -1189 -200 -1177
rect 200 -121 258 -109
rect 200 -1177 212 -121
rect 246 -1177 258 -121
rect 200 -1189 258 -1177
<< ndiffc >>
rect -246 121 -212 1177
rect 212 121 246 1177
rect -246 -1177 -212 -121
rect 212 -1177 246 -121
<< psubdiff >>
rect -360 1329 -264 1363
rect 264 1329 360 1363
rect -360 1267 -326 1329
rect 326 1267 360 1329
rect -360 -1329 -326 -1267
rect 326 -1329 360 -1267
rect -360 -1363 -264 -1329
rect 264 -1363 360 -1329
<< psubdiffcont >>
rect -264 1329 264 1363
rect -360 -1267 -326 1267
rect 326 -1267 360 1267
rect -264 -1363 264 -1329
<< poly >>
rect -200 1261 200 1277
rect -200 1227 -184 1261
rect 184 1227 200 1261
rect -200 1189 200 1227
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -1227 200 -1189
rect -200 -1261 -184 -1227
rect 184 -1261 200 -1227
rect -200 -1277 200 -1261
<< polycont >>
rect -184 1227 184 1261
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -1261 184 -1227
<< locali >>
rect -360 1329 -264 1363
rect 264 1329 360 1363
rect -360 1267 -326 1329
rect 326 1267 360 1329
rect -200 1227 -184 1261
rect 184 1227 200 1261
rect -246 1177 -212 1193
rect -246 105 -212 121
rect 212 1177 246 1193
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -1193 -212 -1177
rect 212 -121 246 -105
rect 212 -1193 246 -1177
rect -200 -1261 -184 -1227
rect 184 -1261 200 -1227
rect -360 -1329 -326 -1267
rect 326 -1329 360 -1267
rect -360 -1363 -264 -1329
rect 264 -1363 360 -1329
<< viali >>
rect -184 1227 184 1261
rect -246 121 -212 1177
rect 212 121 246 1177
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -1177 -212 -121
rect 212 -1177 246 -121
rect -184 -1261 184 -1227
<< metal1 >>
rect -196 1261 196 1267
rect -196 1227 -184 1261
rect 184 1227 196 1261
rect -196 1221 196 1227
rect -252 1177 -206 1189
rect -252 121 -246 1177
rect -212 121 -206 1177
rect -252 109 -206 121
rect 206 1177 252 1189
rect 206 121 212 1177
rect 246 121 252 1177
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -1177 -246 -121
rect -212 -1177 -206 -121
rect -252 -1189 -206 -1177
rect 206 -121 252 -109
rect 206 -1177 212 -121
rect 246 -1177 252 -121
rect 206 -1189 252 -1177
rect -196 -1227 196 -1221
rect -196 -1261 -184 -1227
rect 184 -1261 196 -1227
rect -196 -1267 196 -1261
<< properties >>
string FIXED_BBOX -343 -1346 343 1346
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.4 l 2 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
