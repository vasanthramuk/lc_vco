* SPICE3 file created from trial.ext - technology: sky130A

.subckt trial gnd
X0 gnd curgate curgate gnd sky130_fd_pr__nfet_01v8 ad=2.5752e+13p pd=1.8804e+08u as=0p ps=0u w=5.4e+06u l=1e+06u
X1 gnd curgate curgate gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X2 gnd VDD VDD gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X3 gnd VDD VDD gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X4 VDD VDD gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X5 gnd VDD VDD gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X6 VDD VDD gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X7 gnd VDD VDD gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X8 VDD VDD gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X9 VDD VDD gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X10 VDD vcntrl gnd sky130_fd_pr__cap_var_lvt w=1e+07u l=500000u
X11 VDD vcntrl gnd sky130_fd_pr__cap_var_lvt w=1e+07u l=500000u
X12 VDD VDD sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X13 VDD VDD sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X14 VDD VDD sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X15 VDD VDD sky130_fd_pr__cap_mim_m3_1 l=2.263e+07u w=2.263e+07u
X16 gnd curgate gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X17 gnd curgate gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X18 gnd curgate gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X19 gnd curgate gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X20 gnd curgate gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
C0 VDD curgate 2.19fF
C1 VDD vcntrl 5.46fF
C2 curgate gnd 6.25fF **FLOATING
C3 VDD gnd 63.88fF **FLOATING
C4 vcntrl gnd 9.28fF **FLOATING
.ends
