magic
tech sky130A
magscale 1 2
timestamp 1671093175
<< error_p >>
rect -43 1086 -37 1092
rect 39 1086 45 1092
rect -49 1080 -43 1086
rect 45 1080 51 1086
rect -49 1026 -43 1032
rect 45 1026 51 1032
rect -43 1020 -37 1026
rect 39 1020 45 1026
<< nwell >>
rect -183 -1091 183 1091
<< pwell >>
rect -293 1091 293 1201
rect -293 -1091 -183 1091
rect 183 -1091 293 1091
rect -293 -1201 293 -1091
<< varactor >>
rect -50 -1000 50 1000
<< psubdiff >>
rect -257 1131 -161 1165
rect 161 1131 257 1165
rect -257 1069 -223 1131
rect 223 1069 257 1131
rect -257 -1131 -223 -1069
rect 223 -1131 257 -1069
rect -257 -1165 -161 -1131
rect 161 -1165 257 -1131
<< nsubdiff >>
rect -147 976 -50 1000
rect -147 -976 -135 976
rect -101 -976 -50 976
rect -147 -1000 -50 -976
rect 50 976 147 1000
rect 50 -976 101 976
rect 135 -976 147 976
rect 50 -1000 147 -976
<< psubdiffcont >>
rect -161 1131 161 1165
rect -257 -1069 -223 1069
rect 223 -1069 257 1069
rect -161 -1165 161 -1131
<< nsubdiffcont >>
rect -135 -976 -101 976
rect 101 -976 135 976
<< poly >>
rect -50 1072 50 1088
rect -50 1038 -34 1072
rect 34 1038 50 1072
rect -50 1000 50 1038
rect -50 -1038 50 -1000
rect -50 -1072 -34 -1038
rect 34 -1072 50 -1038
rect -50 -1088 50 -1072
<< polycont >>
rect -34 1038 34 1072
rect -34 -1072 34 -1038
<< locali >>
rect -257 1131 -161 1165
rect 161 1131 257 1165
rect -257 1069 -223 1131
rect -50 1038 -34 1072
rect 34 1038 50 1072
rect 223 1069 257 1131
rect -135 976 -101 992
rect -135 -992 -101 -976
rect 101 976 135 992
rect 101 -992 135 -976
rect -257 -1131 -223 -1069
rect -50 -1072 -34 -1038
rect 34 -1072 50 -1038
rect 223 -1131 257 -1069
rect -257 -1165 -161 -1131
rect 161 -1165 257 -1131
<< viali >>
rect -34 1038 34 1072
rect -135 -976 -101 976
rect 101 -976 135 976
rect -34 -1072 34 -1038
<< metal1 >>
rect -57 1086 61 1092
rect -57 1026 -43 1086
rect 45 1026 61 1086
rect -57 1014 61 1026
rect -141 976 -95 988
rect -141 -976 -135 976
rect -101 -976 -95 976
rect -141 -988 -95 -976
rect 95 976 141 988
rect 95 -976 101 976
rect 135 -976 141 976
rect 95 -988 141 -976
rect -46 -1038 46 -1032
rect -46 -1072 -34 -1038
rect 34 -1072 46 -1038
rect -46 -1078 46 -1072
<< via1 >>
rect -43 1072 45 1086
rect -43 1038 -34 1072
rect -34 1038 34 1072
rect 34 1038 45 1072
rect -43 1026 45 1038
<< properties >>
string FIXED_BBOX -240 -1148 240 1148
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 10 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
