magic
tech sky130A
magscale 1 2
timestamp 1671089082
<< pwell >>
rect -683 -1119 683 1119
<< nmos >>
rect -487 109 -287 909
rect -229 109 -29 909
rect 29 109 229 909
rect 287 109 487 909
rect -487 -909 -287 -109
rect -229 -909 -29 -109
rect 29 -909 229 -109
rect 287 -909 487 -109
<< ndiff >>
rect -545 897 -487 909
rect -545 121 -533 897
rect -499 121 -487 897
rect -545 109 -487 121
rect -287 897 -229 909
rect -287 121 -275 897
rect -241 121 -229 897
rect -287 109 -229 121
rect -29 897 29 909
rect -29 121 -17 897
rect 17 121 29 897
rect -29 109 29 121
rect 229 897 287 909
rect 229 121 241 897
rect 275 121 287 897
rect 229 109 287 121
rect 487 897 545 909
rect 487 121 499 897
rect 533 121 545 897
rect 487 109 545 121
rect -545 -121 -487 -109
rect -545 -897 -533 -121
rect -499 -897 -487 -121
rect -545 -909 -487 -897
rect -287 -121 -229 -109
rect -287 -897 -275 -121
rect -241 -897 -229 -121
rect -287 -909 -229 -897
rect -29 -121 29 -109
rect -29 -897 -17 -121
rect 17 -897 29 -121
rect -29 -909 29 -897
rect 229 -121 287 -109
rect 229 -897 241 -121
rect 275 -897 287 -121
rect 229 -909 287 -897
rect 487 -121 545 -109
rect 487 -897 499 -121
rect 533 -897 545 -121
rect 487 -909 545 -897
<< ndiffc >>
rect -533 121 -499 897
rect -275 121 -241 897
rect -17 121 17 897
rect 241 121 275 897
rect 499 121 533 897
rect -533 -897 -499 -121
rect -275 -897 -241 -121
rect -17 -897 17 -121
rect 241 -897 275 -121
rect 499 -897 533 -121
<< psubdiff >>
rect -647 1049 -551 1083
rect 551 1049 647 1083
rect -647 987 -613 1049
rect 613 987 647 1049
rect -647 -1049 -613 -987
rect 613 -1049 647 -987
rect -647 -1083 -551 -1049
rect 551 -1083 647 -1049
<< psubdiffcont >>
rect -551 1049 551 1083
rect -647 -987 -613 987
rect 613 -987 647 987
rect -551 -1083 551 -1049
<< poly >>
rect -487 981 -287 997
rect -487 947 -471 981
rect -303 947 -287 981
rect -487 909 -287 947
rect -229 981 -29 997
rect -229 947 -213 981
rect -45 947 -29 981
rect -229 909 -29 947
rect 29 981 229 997
rect 29 947 45 981
rect 213 947 229 981
rect 29 909 229 947
rect 287 981 487 997
rect 287 947 303 981
rect 471 947 487 981
rect 287 909 487 947
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect -487 -947 -287 -909
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -487 -997 -287 -981
rect -229 -947 -29 -909
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect -229 -997 -29 -981
rect 29 -947 229 -909
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 29 -997 229 -981
rect 287 -947 487 -909
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 287 -997 487 -981
<< polycont >>
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
<< locali >>
rect -647 1049 -551 1083
rect 551 1049 647 1083
rect -647 987 -613 1049
rect 613 987 647 1049
rect -487 947 -471 981
rect -303 947 -287 981
rect -229 947 -213 981
rect -45 947 -29 981
rect 29 947 45 981
rect 213 947 229 981
rect 287 947 303 981
rect 471 947 487 981
rect -533 897 -499 913
rect -275 897 -241 913
rect -284 360 -275 382
rect -17 897 17 913
rect 241 897 275 913
rect -241 360 -230 382
rect -232 334 -230 360
rect -533 105 -499 121
rect -275 105 -241 121
rect 230 360 241 382
rect 499 897 533 913
rect 275 360 284 382
rect 230 334 232 360
rect -17 105 17 121
rect 241 105 275 121
rect 499 105 533 121
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect -533 -121 -499 -105
rect -275 -121 -241 -105
rect -17 -121 17 -105
rect -533 -913 -499 -897
rect 241 -121 275 -105
rect 499 -121 533 -105
rect -275 -913 -241 -897
rect -17 -913 17 -897
rect 241 -913 275 -897
rect 499 -913 533 -897
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 287 -981 303 -947
rect 471 -981 487 -947
rect -647 -1049 -613 -987
rect 613 -1049 647 -987
rect -647 -1083 -551 -1049
rect 551 -1083 647 -1049
<< viali >>
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect -648 652 -647 822
rect -647 652 -613 822
rect -613 652 -612 822
rect -542 658 -533 824
rect -533 658 -499 824
rect -499 658 -490 824
rect -24 706 -17 822
rect -26 658 -17 706
rect -24 656 -17 658
rect -17 656 17 822
rect 17 656 28 822
rect -284 306 -275 360
rect -275 306 -241 360
rect -241 306 -232 360
rect 492 658 499 824
rect 499 658 533 824
rect 533 658 544 824
rect 232 306 241 360
rect 241 306 275 360
rect 275 306 284 360
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect -280 -380 -275 -318
rect -275 -380 -241 -318
rect -241 -380 -232 -318
rect -540 -828 -533 -660
rect -533 -828 -499 -660
rect -499 -828 -488 -660
rect 234 -378 241 -316
rect 241 -378 275 -316
rect 275 -378 282 -316
rect -26 -820 -17 -666
rect -17 -820 17 -666
rect 17 -820 26 -666
rect 488 -820 499 -666
rect 499 -820 533 -666
rect 533 -820 542 -666
rect 594 -820 613 -666
rect 613 -820 647 -666
rect 647 -820 648 -666
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
<< metal1 >>
rect -296 987 -206 988
rect -38 987 58 988
rect 216 987 310 988
rect -483 981 483 987
rect -483 947 -471 981
rect -303 947 -213 981
rect -45 947 45 981
rect 213 947 303 981
rect 471 947 483 981
rect -483 941 483 947
rect -296 940 -206 941
rect -38 940 58 941
rect 216 940 310 941
rect -666 824 558 836
rect -666 822 -542 824
rect -666 652 -648 822
rect -612 658 -542 822
rect -490 822 492 824
rect -490 706 -24 822
rect -490 658 -26 706
rect 28 658 492 822
rect 544 658 558 824
rect -612 656 -24 658
rect 28 656 558 658
rect -612 652 558 656
rect -666 638 558 652
rect -298 368 -234 380
rect -298 366 306 368
rect -298 360 84 366
rect -298 306 -284 360
rect -232 306 84 360
rect -298 300 84 306
rect 142 360 306 366
rect 142 306 232 360
rect 284 306 306 360
rect 142 300 306 306
rect -298 298 306 300
rect -298 292 -234 298
rect -164 84 -88 102
rect -300 77 -198 78
rect -164 77 -154 84
rect -483 71 -154 77
rect -96 77 -88 84
rect -38 77 54 78
rect 218 77 318 78
rect -96 71 483 77
rect -483 37 -471 71
rect -303 37 -213 71
rect -45 37 45 71
rect 213 37 303 71
rect 471 37 483 71
rect -483 31 -154 37
rect -300 30 -198 31
rect -164 30 -154 31
rect -96 31 483 37
rect -96 30 -88 31
rect -38 30 54 31
rect 218 30 318 31
rect -164 16 -88 30
rect 72 -22 152 -14
rect 72 -30 84 -22
rect -298 -31 -210 -30
rect -42 -31 84 -30
rect -483 -37 84 -31
rect 142 -31 152 -22
rect 214 -31 308 -30
rect 142 -37 483 -31
rect -483 -71 -471 -37
rect -303 -71 -213 -37
rect -45 -71 45 -37
rect 213 -71 303 -37
rect 471 -71 483 -37
rect -483 -77 84 -71
rect -298 -78 -210 -77
rect -42 -78 84 -77
rect 72 -88 84 -78
rect 142 -77 483 -71
rect 142 -88 152 -77
rect 214 -78 308 -77
rect 72 -96 152 -88
rect -294 -308 -238 -300
rect 228 -308 298 -300
rect -294 -316 298 -308
rect -294 -318 234 -316
rect -294 -380 -280 -318
rect -232 -322 234 -318
rect -232 -376 -154 -322
rect -96 -376 234 -322
rect -232 -378 234 -376
rect 282 -378 298 -316
rect -232 -380 298 -378
rect -294 -388 298 -380
rect -294 -394 -238 -388
rect 228 -394 298 -388
rect -556 -660 656 -646
rect -556 -828 -540 -660
rect -488 -666 656 -660
rect -488 -820 -26 -666
rect 26 -820 488 -666
rect 542 -820 594 -666
rect 648 -820 656 -666
rect -488 -828 656 -820
rect -556 -842 656 -828
rect -298 -941 -214 -940
rect -42 -941 44 -940
rect 218 -941 296 -940
rect -483 -947 483 -941
rect -483 -981 -471 -947
rect -303 -981 -213 -947
rect -45 -981 45 -947
rect 213 -981 303 -947
rect 471 -981 483 -947
rect -483 -987 483 -981
rect -298 -988 -214 -987
rect -42 -988 44 -987
rect 218 -988 296 -987
<< via1 >>
rect 84 300 142 366
rect -154 71 -96 84
rect -154 37 -96 71
rect -154 30 -96 37
rect 84 -37 142 -22
rect 84 -71 142 -37
rect 84 -88 142 -71
rect -154 -376 -96 -322
<< metal2 >>
rect 72 366 154 386
rect 72 300 84 366
rect 142 300 154 366
rect -170 84 -86 104
rect -170 30 -154 84
rect -96 30 -86 84
rect -170 -322 -86 30
rect 72 -22 154 300
rect 72 -88 84 -22
rect 142 -88 154 -22
rect 72 -100 154 -88
rect -170 -376 -154 -322
rect -96 -376 -86 -322
rect -170 -390 -86 -376
<< properties >>
string FIXED_BBOX -630 -1066 630 1066
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 1 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
