magic
tech sky130A
magscale 1 2
timestamp 1670750879
<< error_p >>
rect 260 41 371 43
<< pwell >>
rect -296 -3346 296 3346
<< nmos >>
rect -100 2056 100 3136
rect -100 758 100 1838
rect -100 -540 100 540
rect -100 -1838 100 -758
rect -100 -3136 100 -2056
<< ndiff >>
rect -158 3124 -100 3136
rect -158 2068 -146 3124
rect -112 2068 -100 3124
rect -158 2056 -100 2068
rect 100 3124 158 3136
rect 100 2069 112 3124
rect 146 2069 158 3124
rect 100 2056 158 2069
rect -158 1826 -100 1838
rect -158 770 -146 1826
rect -112 770 -100 1826
rect -158 758 -100 770
rect 100 1826 158 1838
rect 100 770 112 1826
rect 146 770 158 1826
rect 100 758 158 770
rect -158 528 -100 540
rect -158 -528 -146 528
rect -112 -528 -100 528
rect -158 -540 -100 -528
rect 100 528 158 540
rect 100 -528 112 528
rect 146 -528 158 528
rect 100 -540 158 -528
rect -158 -770 -100 -758
rect -158 -1826 -146 -770
rect -112 -1826 -100 -770
rect -158 -1838 -100 -1826
rect 100 -770 158 -758
rect 100 -1826 112 -770
rect 146 -1826 158 -770
rect 100 -1838 158 -1826
rect -158 -2068 -100 -2056
rect -158 -3124 -146 -2068
rect -112 -3124 -100 -2068
rect -158 -3136 -100 -3124
rect 100 -2068 158 -2056
rect 100 -3124 112 -2068
rect 146 -3124 158 -2068
rect 100 -3136 158 -3124
<< ndiffc >>
rect -146 2068 -112 3124
rect 112 2069 146 3124
rect -146 770 -112 1826
rect 112 770 146 1826
rect -146 -528 -112 528
rect 112 -528 146 528
rect -146 -1826 -112 -770
rect 112 -1826 146 -770
rect -146 -3124 -112 -2068
rect 112 -3124 146 -2068
<< psubdiff >>
rect -260 3276 -164 3310
rect 164 3276 260 3310
rect -260 3214 -226 3276
rect 226 3214 260 3276
rect -260 -3276 -226 -3214
rect 226 -3276 260 -3214
rect -260 -3310 -164 -3276
rect 164 -3310 260 -3276
<< psubdiffcont >>
rect -164 3276 164 3310
rect -260 -3214 -226 3214
rect 226 -3214 260 3214
rect -164 -3310 164 -3276
<< poly >>
rect -100 3208 100 3224
rect -100 3174 -84 3208
rect 84 3174 100 3208
rect -100 3136 100 3174
rect -100 1968 100 2056
rect -99 1926 99 1968
rect -100 1838 100 1926
rect -100 670 100 758
rect -99 628 99 670
rect -100 540 100 628
rect -100 -628 100 -540
rect -99 -670 99 -628
rect -100 -758 100 -670
rect -100 -1926 100 -1838
rect -99 -1968 99 -1926
rect -100 -2056 100 -1968
rect -100 -3174 100 -3136
rect -100 -3208 -84 -3174
rect 84 -3208 100 -3174
rect -100 -3224 100 -3208
<< polycont >>
rect -84 3174 84 3208
rect -84 -3208 84 -3174
<< locali >>
rect -260 3276 -164 3310
rect 164 3276 260 3310
rect -260 3214 -226 3276
rect 226 3214 260 3276
rect -100 3174 -84 3208
rect 84 3174 100 3208
rect -146 3124 -112 3140
rect 112 3124 146 3140
rect -146 2052 -112 2068
rect 111 2069 112 2073
rect 146 2069 149 2073
rect -146 1826 -112 1842
rect 111 1826 149 2069
rect 111 1825 112 1826
rect -146 754 -112 770
rect 146 1825 149 1826
rect 146 770 147 780
rect -146 528 -112 544
rect -146 -544 -112 -528
rect 112 533 147 770
rect 112 528 146 533
rect 146 9 226 43
rect 112 -537 146 -528
rect -146 -770 -112 -754
rect -146 -1842 -112 -1826
rect 112 -759 149 -537
rect 112 -770 146 -759
rect 146 -1826 152 -1808
rect 112 -1842 152 -1826
rect 113 -2052 152 -1842
rect -146 -2068 -112 -2052
rect -146 -3140 -112 -3124
rect 112 -2062 152 -2052
rect 112 -2065 149 -2062
rect 112 -2068 146 -2065
rect 112 -3140 146 -3124
rect -100 -3208 -84 -3174
rect 84 -3208 100 -3174
rect -260 -3276 -226 -3214
rect 260 9 371 41
rect 226 -3276 260 -3214
rect -260 -3310 -164 -3276
rect 164 -3310 260 -3276
<< viali >>
rect -146 2068 -112 3124
rect -146 770 -112 1826
rect -146 -528 -112 528
rect -146 -1826 -112 -770
rect -146 -2719 -112 -2068
rect -84 -3208 84 -3174
<< metal1 >>
rect -157 3125 -99 3165
rect -157 3124 -101 3125
rect -157 2068 -146 3124
rect -112 2068 -101 3124
rect -157 2055 -101 2068
rect -146 1849 -110 2055
rect -163 1826 -99 1849
rect -163 1809 -146 1826
rect -157 770 -146 1809
rect -112 1809 -99 1826
rect -112 770 -101 1809
rect -157 755 -101 770
rect -157 543 -114 755
rect -157 528 -101 543
rect -157 25 -146 528
rect -449 -25 -146 25
rect -157 -513 -146 -25
rect -159 -528 -146 -513
rect -112 -513 -101 528
rect -112 -528 -99 -513
rect -159 -559 -99 -528
rect -144 -757 -113 -559
rect -157 -770 -99 -757
rect -157 -1826 -146 -770
rect -112 -1826 -99 -770
rect -157 -1841 -99 -1826
rect -157 -2055 -128 -1841
rect -159 -2068 -103 -2055
rect -159 -2719 -146 -2068
rect -112 -2719 -103 -2068
rect -157 -2761 -103 -2719
rect -99 -3174 99 -3159
rect -99 -3208 -84 -3174
rect 84 -3208 99 -3174
rect -99 -3225 99 -3208
rect -29 -3571 15 -3225
<< labels >>
rlabel metal1 -441 -17 -415 23 1 vp
rlabel locali 359 11 369 35 1 gnd
rlabel metal1 -19 -3563 5 -3539 1 cursrc1gate
<< properties >>
string FIXED_BBOX -243 -3293 243 3293
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.4 l 1 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
