magic
tech sky130A
magscale 1 2
timestamp 1671513803
<< error_p >>
rect -87 3210 91 3216
rect -87 3181 -81 3210
rect 85 3181 91 3210
rect -87 3175 91 3181
<< pwell >>
rect -296 -3346 296 3346
<< nmos >>
rect -100 2056 100 3136
rect -100 758 100 1838
rect -100 -540 100 540
rect -100 -1838 100 -758
rect -100 -3136 100 -2056
<< ndiff >>
rect -158 3124 -100 3136
rect -158 2068 -146 3124
rect -112 2068 -100 3124
rect -158 2056 -100 2068
rect 100 3124 158 3136
rect 100 2068 112 3124
rect 146 2068 158 3124
rect 100 2056 158 2068
rect -158 1826 -100 1838
rect -158 770 -146 1826
rect -112 770 -100 1826
rect -158 758 -100 770
rect 100 1826 158 1838
rect 100 770 112 1826
rect 146 770 158 1826
rect 100 758 158 770
rect -158 528 -100 540
rect -158 -528 -146 528
rect -112 -528 -100 528
rect -158 -540 -100 -528
rect 100 528 158 540
rect 100 -528 112 528
rect 146 -528 158 528
rect 100 -540 158 -528
rect -158 -770 -100 -758
rect -158 -1826 -146 -770
rect -112 -1826 -100 -770
rect -158 -1838 -100 -1826
rect 100 -770 158 -758
rect 100 -1826 112 -770
rect 146 -1826 158 -770
rect 100 -1838 158 -1826
rect -158 -2068 -100 -2056
rect -158 -3124 -146 -2068
rect -112 -3124 -100 -2068
rect -158 -3136 -100 -3124
rect 100 -2068 158 -2056
rect 100 -3124 112 -2068
rect 146 -3124 158 -2068
rect 100 -3136 158 -3124
<< ndiffc >>
rect -146 2068 -112 3124
rect 112 2068 146 3124
rect -146 770 -112 1826
rect 112 770 146 1826
rect -146 -528 -112 528
rect 112 -528 146 528
rect -146 -1826 -112 -770
rect 112 -1826 146 -770
rect -146 -3124 -112 -2068
rect 112 -3124 146 -2068
<< psubdiff >>
rect -260 3276 -164 3310
rect 164 3276 260 3310
rect -260 3214 -226 3276
rect 226 3214 260 3276
rect -260 -3276 -226 -3214
rect 226 -3276 260 -3214
rect -260 -3310 -164 -3276
rect 164 -3310 260 -3276
<< psubdiffcont >>
rect -164 3276 164 3310
rect -260 -3214 -226 3214
rect 226 -3214 260 3214
rect -164 -3310 164 -3276
<< poly >>
rect -100 3214 100 3224
rect -100 3179 -84 3214
rect 84 3179 100 3214
rect -100 3136 100 3179
rect -100 1838 100 2056
rect -100 540 100 758
rect -100 -758 100 -540
rect -100 -2056 100 -1838
rect -100 -3224 100 -3136
<< polycont >>
rect -84 3179 84 3214
<< locali >>
rect -260 3276 -164 3310
rect 164 3276 260 3310
rect -260 3214 -226 3276
rect -100 3216 101 3218
rect -100 3175 -87 3216
rect 91 3175 101 3216
rect -100 3174 101 3175
rect 226 3214 260 3276
rect -146 3124 -112 3140
rect -146 1826 -112 2068
rect -146 528 -112 770
rect -146 -770 -112 -528
rect -146 -2068 -112 -1826
rect -146 -3140 -112 -3124
rect 112 3124 146 3140
rect 112 1826 146 2068
rect 112 528 146 770
rect 112 -770 146 -528
rect 112 -2068 146 -1826
rect 112 -3140 146 -3124
rect -260 -3276 -226 -3214
rect 226 -3276 260 -3214
rect -260 -3310 -164 -3276
rect 164 -3310 260 -3276
<< viali >>
rect -87 3214 91 3216
rect -87 3179 -84 3214
rect -84 3179 84 3214
rect 84 3179 91 3214
rect -87 3175 91 3179
<< properties >>
string FIXED_BBOX -243 -3293 243 3293
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.4 l 1 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
