magic
tech sky130A
magscale 1 2
timestamp 1670046431
<< nwell >>
rect -223 -1131 223 1131
<< pwell >>
rect -514 1131 514 1422
rect -514 -1131 -223 1131
rect 223 -1131 514 1131
rect -514 -1422 514 -1131
<< mvvaractor >>
rect -50 -1000 50 1000
<< mvpsubdiff >>
rect -438 1334 438 1346
rect -438 1300 -330 1334
rect 330 1300 438 1334
rect -438 1288 438 1300
rect -438 1238 -380 1288
rect -438 -1238 -426 1238
rect -392 -1238 -380 1238
rect 380 1238 438 1288
rect -438 -1288 -380 -1238
rect 380 -1238 392 1238
rect 426 -1238 438 1238
rect 380 -1288 438 -1238
rect -438 -1300 438 -1288
rect -438 -1334 -330 -1300
rect 330 -1334 438 -1300
rect -438 -1346 438 -1334
<< mvnsubdiff >>
rect -147 976 -50 1000
rect -147 -976 -135 976
rect -101 -976 -50 976
rect -147 -1000 -50 -976
rect 50 976 147 1000
rect 50 -976 101 976
rect 135 -976 147 976
rect 50 -1000 147 -976
<< mvpsubdiffcont >>
rect -330 1300 330 1334
rect -426 -1238 -392 1238
rect 392 -1238 426 1238
rect -330 -1334 330 -1300
<< mvnsubdiffcont >>
rect -135 -976 -101 976
rect 101 -976 135 976
<< poly >>
rect -50 1072 50 1088
rect -50 1038 -34 1072
rect 34 1038 50 1072
rect -50 1000 50 1038
rect -50 -1038 50 -1000
rect -50 -1072 -34 -1038
rect 34 -1072 50 -1038
rect -50 -1088 50 -1072
<< polycont >>
rect -34 1038 34 1072
rect -34 -1072 34 -1038
<< locali >>
rect -426 1300 -330 1334
rect 330 1300 426 1334
rect -426 1238 -392 1300
rect 392 1238 426 1300
rect -50 1038 -34 1072
rect 34 1038 50 1072
rect -135 976 -101 992
rect -135 -992 -101 -976
rect 101 976 135 992
rect 101 -992 135 -976
rect -50 -1072 -34 -1038
rect 34 -1072 50 -1038
rect -426 -1300 -392 -1238
rect 392 -1300 426 -1238
rect -426 -1334 -330 -1300
rect 330 -1334 426 -1300
<< viali >>
rect -34 1038 34 1072
rect -135 -976 -101 976
rect 101 -976 135 976
rect -34 -1072 34 -1038
<< metal1 >>
rect -46 1072 46 1078
rect -46 1038 -34 1072
rect 34 1038 46 1072
rect -46 1032 46 1038
rect -141 976 -95 988
rect -141 -976 -135 976
rect -101 -976 -95 976
rect -141 -988 -95 -976
rect 95 976 141 988
rect 95 -976 101 976
rect 135 -976 141 976
rect 95 -988 141 -976
rect -46 -1038 46 -1032
rect -46 -1072 -34 -1038
rect 34 -1072 46 -1038
rect -46 -1078 46 -1072
<< properties >>
string FIXED_BBOX -409 -1317 409 1317
string gencell sky130_fd_pr__cap_var
string library sky130
string parameters w 10 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
