magic
tech sky130A
magscale 1 2
timestamp 1670833676
<< nwell >>
rect -2973 -191 -2607 191
rect -2353 -191 -1987 191
rect -1733 -191 -1367 191
rect -1113 -191 -747 191
rect -493 -191 -127 191
rect 127 -191 493 191
rect 747 -191 1113 191
rect 1367 -191 1733 191
rect 1987 -191 2353 191
rect 2607 -191 2973 191
<< pwell >>
rect -3083 191 3083 301
rect -3083 -191 -2973 191
rect -2607 -191 -2353 191
rect -1987 -191 -1733 191
rect -1367 -191 -1113 191
rect -747 -191 -493 191
rect -127 -191 127 191
rect 493 -191 747 191
rect 1113 -191 1367 191
rect 1733 -191 1987 191
rect 2353 -191 2607 191
rect 2973 -191 3083 191
rect -3083 -301 3083 -191
<< varactor >>
rect -2840 -100 -2740 100
rect -2220 -100 -2120 100
rect -1600 -100 -1500 100
rect -980 -100 -880 100
rect -360 -100 -260 100
rect 260 -100 360 100
rect 880 -100 980 100
rect 1500 -100 1600 100
rect 2120 -100 2220 100
rect 2740 -100 2840 100
<< psubdiff >>
rect -3047 231 -2951 265
rect 2951 231 3047 265
rect -3047 169 -3013 231
rect 3013 169 3047 231
rect -3047 -231 -3013 -169
rect 3013 -231 3047 -169
rect -3047 -265 -2951 -231
rect 2951 -265 3047 -231
<< nsubdiff >>
rect -2937 76 -2840 100
rect -2937 -76 -2925 76
rect -2891 -76 -2840 76
rect -2937 -100 -2840 -76
rect -2740 76 -2643 100
rect -2740 -76 -2689 76
rect -2655 -76 -2643 76
rect -2740 -100 -2643 -76
rect -2317 76 -2220 100
rect -2317 -76 -2305 76
rect -2271 -76 -2220 76
rect -2317 -100 -2220 -76
rect -2120 76 -2023 100
rect -2120 -76 -2069 76
rect -2035 -76 -2023 76
rect -2120 -100 -2023 -76
rect -1697 76 -1600 100
rect -1697 -76 -1685 76
rect -1651 -76 -1600 76
rect -1697 -100 -1600 -76
rect -1500 76 -1403 100
rect -1500 -76 -1449 76
rect -1415 -76 -1403 76
rect -1500 -100 -1403 -76
rect -1077 76 -980 100
rect -1077 -76 -1065 76
rect -1031 -76 -980 76
rect -1077 -100 -980 -76
rect -880 76 -783 100
rect -880 -76 -829 76
rect -795 -76 -783 76
rect -880 -100 -783 -76
rect -457 76 -360 100
rect -457 -76 -445 76
rect -411 -76 -360 76
rect -457 -100 -360 -76
rect -260 76 -163 100
rect -260 -76 -209 76
rect -175 -76 -163 76
rect -260 -100 -163 -76
rect 163 76 260 100
rect 163 -76 175 76
rect 209 -76 260 76
rect 163 -100 260 -76
rect 360 76 457 100
rect 360 -76 411 76
rect 445 -76 457 76
rect 360 -100 457 -76
rect 783 76 880 100
rect 783 -76 795 76
rect 829 -76 880 76
rect 783 -100 880 -76
rect 980 76 1077 100
rect 980 -76 1031 76
rect 1065 -76 1077 76
rect 980 -100 1077 -76
rect 1403 76 1500 100
rect 1403 -76 1415 76
rect 1449 -76 1500 76
rect 1403 -100 1500 -76
rect 1600 76 1697 100
rect 1600 -76 1651 76
rect 1685 -76 1697 76
rect 1600 -100 1697 -76
rect 2023 76 2120 100
rect 2023 -76 2035 76
rect 2069 -76 2120 76
rect 2023 -100 2120 -76
rect 2220 76 2317 100
rect 2220 -76 2271 76
rect 2305 -76 2317 76
rect 2220 -100 2317 -76
rect 2643 76 2740 100
rect 2643 -76 2655 76
rect 2689 -76 2740 76
rect 2643 -100 2740 -76
rect 2840 76 2937 100
rect 2840 -76 2891 76
rect 2925 -76 2937 76
rect 2840 -100 2937 -76
<< psubdiffcont >>
rect -2951 231 2951 265
rect -3047 -169 -3013 169
rect 3013 -169 3047 169
rect -2951 -265 2951 -231
<< nsubdiffcont >>
rect -2925 -76 -2891 76
rect -2689 -76 -2655 76
rect -2305 -76 -2271 76
rect -2069 -76 -2035 76
rect -1685 -76 -1651 76
rect -1449 -76 -1415 76
rect -1065 -76 -1031 76
rect -829 -76 -795 76
rect -445 -76 -411 76
rect -209 -76 -175 76
rect 175 -76 209 76
rect 411 -76 445 76
rect 795 -76 829 76
rect 1031 -76 1065 76
rect 1415 -76 1449 76
rect 1651 -76 1685 76
rect 2035 -76 2069 76
rect 2271 -76 2305 76
rect 2655 -76 2689 76
rect 2891 -76 2925 76
<< poly >>
rect -2840 172 -2740 188
rect -2840 138 -2824 172
rect -2756 138 -2740 172
rect -2840 100 -2740 138
rect -2220 172 -2120 188
rect -2220 138 -2204 172
rect -2136 138 -2120 172
rect -2220 100 -2120 138
rect -1600 172 -1500 188
rect -1600 138 -1584 172
rect -1516 138 -1500 172
rect -1600 100 -1500 138
rect -980 172 -880 188
rect -980 138 -964 172
rect -896 138 -880 172
rect -980 100 -880 138
rect -360 172 -260 188
rect -360 138 -344 172
rect -276 138 -260 172
rect -360 100 -260 138
rect 260 172 360 188
rect 260 138 276 172
rect 344 138 360 172
rect 260 100 360 138
rect 880 172 980 188
rect 880 138 896 172
rect 964 138 980 172
rect 880 100 980 138
rect 1500 172 1600 188
rect 1500 138 1516 172
rect 1584 138 1600 172
rect 1500 100 1600 138
rect 2120 172 2220 188
rect 2120 138 2136 172
rect 2204 138 2220 172
rect 2120 100 2220 138
rect 2740 172 2840 188
rect 2740 138 2756 172
rect 2824 138 2840 172
rect 2740 100 2840 138
rect -2840 -138 -2740 -100
rect -2840 -172 -2824 -138
rect -2756 -172 -2740 -138
rect -2840 -188 -2740 -172
rect -2220 -138 -2120 -100
rect -2220 -172 -2204 -138
rect -2136 -172 -2120 -138
rect -2220 -188 -2120 -172
rect -1600 -138 -1500 -100
rect -1600 -172 -1584 -138
rect -1516 -172 -1500 -138
rect -1600 -188 -1500 -172
rect -980 -138 -880 -100
rect -980 -172 -964 -138
rect -896 -172 -880 -138
rect -980 -188 -880 -172
rect -360 -138 -260 -100
rect -360 -172 -344 -138
rect -276 -172 -260 -138
rect -360 -188 -260 -172
rect 260 -138 360 -100
rect 260 -172 276 -138
rect 344 -172 360 -138
rect 260 -188 360 -172
rect 880 -138 980 -100
rect 880 -172 896 -138
rect 964 -172 980 -138
rect 880 -188 980 -172
rect 1500 -138 1600 -100
rect 1500 -172 1516 -138
rect 1584 -172 1600 -138
rect 1500 -188 1600 -172
rect 2120 -138 2220 -100
rect 2120 -172 2136 -138
rect 2204 -172 2220 -138
rect 2120 -188 2220 -172
rect 2740 -138 2840 -100
rect 2740 -172 2756 -138
rect 2824 -172 2840 -138
rect 2740 -188 2840 -172
<< polycont >>
rect -2824 138 -2756 172
rect -2204 138 -2136 172
rect -1584 138 -1516 172
rect -964 138 -896 172
rect -344 138 -276 172
rect 276 138 344 172
rect 896 138 964 172
rect 1516 138 1584 172
rect 2136 138 2204 172
rect 2756 138 2824 172
rect -2824 -172 -2756 -138
rect -2204 -172 -2136 -138
rect -1584 -172 -1516 -138
rect -964 -172 -896 -138
rect -344 -172 -276 -138
rect 276 -172 344 -138
rect 896 -172 964 -138
rect 1516 -172 1584 -138
rect 2136 -172 2204 -138
rect 2756 -172 2824 -138
<< locali >>
rect -3047 231 -2951 265
rect 2951 231 3047 265
rect -3047 169 -3013 231
rect -2840 138 -2824 172
rect -2756 138 -2740 172
rect -2220 138 -2204 172
rect -2136 138 -2120 172
rect -1600 138 -1584 172
rect -1516 138 -1500 172
rect -980 138 -964 172
rect -896 138 -880 172
rect -360 138 -344 172
rect -276 138 -260 172
rect 260 138 276 172
rect 344 138 360 172
rect 880 138 896 172
rect 964 138 980 172
rect 1500 138 1516 172
rect 1584 138 1600 172
rect 2120 138 2136 172
rect 2204 138 2220 172
rect 2740 138 2756 172
rect 2824 138 2840 172
rect 3013 169 3047 231
rect -2925 76 -2891 92
rect -2925 -92 -2891 -76
rect -2689 76 -2655 92
rect -2689 -92 -2655 -76
rect -2305 76 -2271 92
rect -2305 -92 -2271 -76
rect -2069 76 -2035 92
rect -2069 -92 -2035 -76
rect -1685 76 -1651 92
rect -1685 -92 -1651 -76
rect -1449 76 -1415 92
rect -1449 -92 -1415 -76
rect -1065 76 -1031 92
rect -1065 -92 -1031 -76
rect -829 76 -795 92
rect -829 -92 -795 -76
rect -445 76 -411 92
rect -445 -92 -411 -76
rect -209 76 -175 92
rect -209 -92 -175 -76
rect 175 76 209 92
rect 175 -92 209 -76
rect 411 76 445 92
rect 411 -92 445 -76
rect 795 76 829 92
rect 795 -92 829 -76
rect 1031 76 1065 92
rect 1031 -92 1065 -76
rect 1415 76 1449 92
rect 1415 -92 1449 -76
rect 1651 76 1685 92
rect 1651 -92 1685 -76
rect 2035 76 2069 92
rect 2035 -92 2069 -76
rect 2271 76 2305 92
rect 2271 -92 2305 -76
rect 2655 76 2689 92
rect 2655 -92 2689 -76
rect 2891 76 2925 92
rect 2891 -92 2925 -76
rect -3047 -231 -3013 -169
rect -2840 -172 -2824 -138
rect -2756 -172 -2740 -138
rect -2220 -172 -2204 -138
rect -2136 -172 -2120 -138
rect -1600 -172 -1584 -138
rect -1516 -172 -1500 -138
rect -980 -172 -964 -138
rect -896 -172 -880 -138
rect -360 -172 -344 -138
rect -276 -172 -260 -138
rect 260 -172 276 -138
rect 344 -172 360 -138
rect 880 -172 896 -138
rect 964 -172 980 -138
rect 1500 -172 1516 -138
rect 1584 -172 1600 -138
rect 2120 -172 2136 -138
rect 2204 -172 2220 -138
rect 2740 -172 2756 -138
rect 2824 -172 2840 -138
rect 3013 -231 3047 -169
rect -3047 -265 -2951 -231
rect 2951 -265 3047 -231
<< viali >>
rect -2824 138 -2756 172
rect -2204 138 -2136 172
rect -1584 138 -1516 172
rect -964 138 -896 172
rect -344 138 -276 172
rect 276 138 344 172
rect 896 138 964 172
rect 1516 138 1584 172
rect 2136 138 2204 172
rect 2756 138 2824 172
rect -2925 -76 -2891 76
rect -2689 -76 -2655 76
rect -2305 -76 -2271 76
rect -2069 -76 -2035 76
rect -1685 -76 -1651 76
rect -1449 -76 -1415 76
rect -1065 -76 -1031 76
rect -829 -76 -795 76
rect -445 -76 -411 76
rect -209 -76 -175 76
rect 175 -76 209 76
rect 411 -76 445 76
rect 795 -76 829 76
rect 1031 -76 1065 76
rect 1415 -76 1449 76
rect 1651 -76 1685 76
rect 2035 -76 2069 76
rect 2271 -76 2305 76
rect 2655 -76 2689 76
rect 2891 -76 2925 76
rect -2824 -172 -2756 -138
rect -2204 -172 -2136 -138
rect -1584 -172 -1516 -138
rect -964 -172 -896 -138
rect -344 -172 -276 -138
rect 276 -172 344 -138
rect 896 -172 964 -138
rect 1516 -172 1584 -138
rect 2136 -172 2204 -138
rect 2756 -172 2824 -138
<< metal1 >>
rect -2836 172 -2744 178
rect -2836 138 -2824 172
rect -2756 138 -2744 172
rect -2836 132 -2744 138
rect -2216 172 -2124 178
rect -2216 138 -2204 172
rect -2136 138 -2124 172
rect -2216 132 -2124 138
rect -1596 172 -1504 178
rect -1596 138 -1584 172
rect -1516 138 -1504 172
rect -1596 132 -1504 138
rect -976 172 -884 178
rect -976 138 -964 172
rect -896 138 -884 172
rect -976 132 -884 138
rect -356 172 -264 178
rect -356 138 -344 172
rect -276 138 -264 172
rect -356 132 -264 138
rect 264 172 356 178
rect 264 138 276 172
rect 344 138 356 172
rect 264 132 356 138
rect 884 172 976 178
rect 884 138 896 172
rect 964 138 976 172
rect 884 132 976 138
rect 1504 172 1596 178
rect 1504 138 1516 172
rect 1584 138 1596 172
rect 1504 132 1596 138
rect 2124 172 2216 178
rect 2124 138 2136 172
rect 2204 138 2216 172
rect 2124 132 2216 138
rect 2744 172 2836 178
rect 2744 138 2756 172
rect 2824 138 2836 172
rect 2744 132 2836 138
rect -2931 76 -2885 88
rect -2931 -76 -2925 76
rect -2891 -76 -2885 76
rect -2931 -88 -2885 -76
rect -2695 76 -2649 88
rect -2695 -76 -2689 76
rect -2655 -76 -2649 76
rect -2695 -88 -2649 -76
rect -2311 76 -2265 88
rect -2311 -76 -2305 76
rect -2271 -76 -2265 76
rect -2311 -88 -2265 -76
rect -2075 76 -2029 88
rect -2075 -76 -2069 76
rect -2035 -76 -2029 76
rect -2075 -88 -2029 -76
rect -1691 76 -1645 88
rect -1691 -76 -1685 76
rect -1651 -76 -1645 76
rect -1691 -88 -1645 -76
rect -1455 76 -1409 88
rect -1455 -76 -1449 76
rect -1415 -76 -1409 76
rect -1455 -88 -1409 -76
rect -1071 76 -1025 88
rect -1071 -76 -1065 76
rect -1031 -76 -1025 76
rect -1071 -88 -1025 -76
rect -835 76 -789 88
rect -835 -76 -829 76
rect -795 -76 -789 76
rect -835 -88 -789 -76
rect -451 76 -405 88
rect -451 -76 -445 76
rect -411 -76 -405 76
rect -451 -88 -405 -76
rect -215 76 -169 88
rect -215 -76 -209 76
rect -175 -76 -169 76
rect -215 -88 -169 -76
rect 169 76 215 88
rect 169 -76 175 76
rect 209 -76 215 76
rect 169 -88 215 -76
rect 405 76 451 88
rect 405 -76 411 76
rect 445 -76 451 76
rect 405 -88 451 -76
rect 789 76 835 88
rect 789 -76 795 76
rect 829 -76 835 76
rect 789 -88 835 -76
rect 1025 76 1071 88
rect 1025 -76 1031 76
rect 1065 -76 1071 76
rect 1025 -88 1071 -76
rect 1409 76 1455 88
rect 1409 -76 1415 76
rect 1449 -76 1455 76
rect 1409 -88 1455 -76
rect 1645 76 1691 88
rect 1645 -76 1651 76
rect 1685 -76 1691 76
rect 1645 -88 1691 -76
rect 2029 76 2075 88
rect 2029 -76 2035 76
rect 2069 -76 2075 76
rect 2029 -88 2075 -76
rect 2265 76 2311 88
rect 2265 -76 2271 76
rect 2305 -76 2311 76
rect 2265 -88 2311 -76
rect 2649 76 2695 88
rect 2649 -76 2655 76
rect 2689 -76 2695 76
rect 2649 -88 2695 -76
rect 2885 76 2931 88
rect 2885 -76 2891 76
rect 2925 -76 2931 76
rect 2885 -88 2931 -76
rect -2836 -138 -2744 -132
rect -2836 -172 -2824 -138
rect -2756 -172 -2744 -138
rect -2836 -178 -2744 -172
rect -2216 -138 -2124 -132
rect -2216 -172 -2204 -138
rect -2136 -172 -2124 -138
rect -2216 -178 -2124 -172
rect -1596 -138 -1504 -132
rect -1596 -172 -1584 -138
rect -1516 -172 -1504 -138
rect -1596 -178 -1504 -172
rect -976 -138 -884 -132
rect -976 -172 -964 -138
rect -896 -172 -884 -138
rect -976 -178 -884 -172
rect -356 -138 -264 -132
rect -356 -172 -344 -138
rect -276 -172 -264 -138
rect -356 -178 -264 -172
rect 264 -138 356 -132
rect 264 -172 276 -138
rect 344 -172 356 -138
rect 264 -178 356 -172
rect 884 -138 976 -132
rect 884 -172 896 -138
rect 964 -172 976 -138
rect 884 -178 976 -172
rect 1504 -138 1596 -132
rect 1504 -172 1516 -138
rect 1584 -172 1596 -138
rect 1504 -178 1596 -172
rect 2124 -138 2216 -132
rect 2124 -172 2136 -138
rect 2204 -172 2216 -138
rect 2124 -178 2216 -172
rect 2744 -138 2836 -132
rect 2744 -172 2756 -138
rect 2824 -172 2836 -138
rect 2744 -178 2836 -172
<< properties >>
string FIXED_BBOX -3030 -248 3030 248
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 1.0 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
