* SPICE3 file created from trial.ext - technology: sky130A

X0 gnd curgate curgate gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X1 gnd curgate curgate gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X2 gnd curgate vp gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X3 gnd curgate vp gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X4 gnd curgate vp gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X5 gnd curgate vp gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
X6 gnd curgate vp gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=1e+06u
C0 vp gnd 5.03fF **FLOATING
C1 curgate gnd 5.68fF **FLOATING
