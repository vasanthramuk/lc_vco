** sch_path: /home/luminatrix/Documents/designs/lc_vco/final.sch
**.subckt final
XC5 vout_m vcntrl GND sky130_fd_pr__cap_var_lvt W=10 L=0.5 VM=1 m=1
XC6 vout_p vcntrl GND sky130_fd_pr__cap_var_lvt W=10 L=0.5 VM=1 m=1
XM1 vout_p vout_m vp vp sky130_fd_pr__nfet_01v8 L=1 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vout_m vout_p vp vp sky130_fd_pr__nfet_01v8 L=1 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1 VDD vout_m sky130_fd_pr__cap_mim_m3_1 W=32 L=32 MF=1 m=1
XC2 VDD vout_p sky130_fd_pr__cap_mim_m3_1 W=32 L=32 MF=1 m=1
XL14 vout_p vout_m VDD GND sky130_fd_pr__ind_05_220
XM3 vp curgate GND GND sky130_fd_pr__nfet_01v8 L=1 W=27 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 idealcs idealcs GND GND sky130_fd_pr__nfet_01v8 L=1 W=10.8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
